BZh91AY&SY޵w ��߀pp��b� ����ak� (����T"�JHziQ@)E*�"���R��(��I)"���(/ 9T

 �"D 
$*!@ ���J�� @ �@�J�   $���� �G    �( �@
 ���}�#���dpz ��K�zԹ�,T�� ���� l�| ��EY���8 �U14���*�P��MS�}�B����iTͽ8��}    >� @  
�(��� �}5�����yiO\��n ������1w4�dWs�]�0��@u*��cc��o0����8 ���!�2轻�����=}��\�}z_|��˞Ξ[�e\ ���    �(e� �=���{�{3�Ҿ۞��� ���˺ڷ9�lq�u�̣ �9o{r^{ z�`���� ����t�{����7��� ���a����\Z�NAǀ�|    �I@Q�� }�I��7<�绔90=���
��@����X>V{p7z ���0�8����Eɡy�>�:w�J���brǽǏj\۞����Jd2[��w;�����^ }�R�  $ ���닮1�s����Q� �c��ϡ�\�rһ��z� �\���Zq��  7��u�y��<�  �������\`�� �z79�>�������q.=        ?H��iT�� �   =IR�  @��E?�U)   LL  �&=��(�*�� �  �O��Cj�U�@� A�� �!T�M52�SLF� =!��'���������_��p���G^���@**���� U] �*���TU_����@�EU���TU]_��R*�����J�*���~r�������7VsP�%�� ����5�&�*�H�#���ö��3[��&MD��a���F��p2|Á�Ԇd&��9������Ì`j"�?�=�y�`�����ro!��	���1��ve��K��s�A�����S)]	��$j���]�M�xk�K�䘙8����5	ܺwbNFꓳVa�a��G�Ύy٭�\�	:�i�8S8��P�7�B��T�h�E�:]�@d��pǇ���[�f(�l۳9ѣ"MNw:09�4�9��I�PƊ����JR��]VW�Ik�&{qs9{i���dMB�
�X�K�X:P���u����
�h�W�n��g�ڞ�|�嫸�*�3�.��[j��ԉ6j"ǣVAPcNF�2m��bh�ib#2q��Şl���TQ�Ć8����Du)B5"Ca��9}�jaڭWH���@�AOR��>)�>g9��\��5�A��޲����d��@��e�uv���D�R���E԰���r�� ��{�0�mקEі�b��#��Պ�*@�)v�c�q(��
�4��SێM�+)A$ÔS���:�@\��J2dc�:�c#-Sj���ģF�`rr1��&��*�AA&��LjN�����KN��;���Y�2p#4=�.A��FX�.��w���)8����GQ8�r{H�0�y��8O���.זv�Ӊ�|�vt��{k"�y��ūP��E{��:���;���V��N'�M�X�T��z�F�v�y�n6���"c'#
�x%	�%	��(J8�ng�h��*�f`m�7	�Ǻuaw�M��n�!�dM�xs����9��Q�r����M���2N�����A���S+H��qȑS׶��P�k|>��y|h~ȋ)�'VRM�4�ۤ�
�����P�e��n)1�L�j-�g3�|�uN4>E+�e��R=�I�,L��|W喊�)@���䆼�����ӳ�ב�;�!(rwY	BP�%	����,��dt���:<6�.��;Xˬ�L���W����U�!���12M����u��bʖ%�	?1,�k�9����R�$�����N�L��3�۫4���v\`	Z�4Re�'�K�Yܮ��sք�n�.��}�U֒kX��%	��%!�G�>�^sN���$"���V����d���K��/P�)
/4�"��;��~�E�;|��c	@h��ƽ�	�L�Xh�:���0�9�"�������;�]��Kr(���5�S�Y]X�tV�p��HN즔u&&N$w`q3\I�,;u8��ٹ���z��05���X�ADC�:���7�b7���.��E���,Ō�Id�L���r�ޞ��哨���.p���\X�!�(�;L�Ȍw��q�)<c-p:á����塋-�NHk7գm���	�d(K�)U�T�R�8���׆�ފ�:�L�&L5ks��tXaĜ'F�sFНBf�6��;��I���q�ƫ�jR!(R�AQA����ջ�}���`ua����z�2WLN�)uN��]/vJ�ti�(���;��˹�9�7��/�Nޓ�d��V@YE�u�Z�Z%a�������A��ŋ[�b��Z�Q*�$���(	P�K�̌-��v..٘�޹���~�D<Y�\Bu��x�/	��i,��tE'vm�a�uΞ�L�u�<�_u<|#Tr��C�I��N��r\7L9ayD����X��%�i��P�6�I�	�%�E,]��h�+4%	T��e�(~Z��v?Y�}:!%�Ԅ��3 �n�Rk05`j���9�x���U�ꮙK)2��K+��3$���RF�[5Iט�r]����NF��ގ�q3������c�[���G��e�c�}���8
�k���*e&T�����N�.�������N��Q��'Y�x��l��\̺��Vt�yk�P�X�'�2P�m���J�J��J����B���j�љ��ѹ�q#''=��>���7'Sdɐj�����a�N�::�g3o.ġ)%�m.Pbi6d%��z��Ց&�y��������p]�b�
�_�"����f�bː��Ժ��[!*����1:��0 �A�H�T�'kS+R$$�E��	N�B4:��[��Дg!��#A���٬t�r1��1+D0ڧP��E��pYŔ���N��
U �����(O3��d%!�!�`fhJ%�6�`�%�!+N�d'P���V�I��WJ	Z�j\�qs{iZ�[^�d�2��͘C�Y���	����N(��J�.�*%��j�/E�E��V�C���<f^^3��л�Y̴�!�a�H�.�JG2�Hs��}My&Γ�L��M�:\��������9����|���k�ѩ�A��G�i�o9	BZ�'#0J�(��O9����٬Ȫwdlt�A��1�&@uff�u	K�'r���b�SW�)�����ђ�A$�k�5	X�BP�%��Q��|㪅���V���V�S<�k#NMڟ�������G`d%`�ԛ��]u�N)����BtP:�H�q��1�a�������:���ׄt43�N�K�g]��њ޸9��N�(��'p��f��2c$�d��GFޖ*�j�ˏ@R��P���b�����SN	9��%x��b�j�j�׺�PbM]����XR�}�L��qv��R�F�i�*_����ܨ�z� ݭ�Z���8�c�5�hrG~^Vv��1V�ި�bVS�f�����Ԅ���6٣|��}
�u�ڜ*�t����Z"cV��U�
K��,C��Os6Q#� �.�)ГI2��{oWEBik�&V͞�ܜL��Ѿm9a��1��:� ��*�zӨ��[�]t�䲔4�������&�K�ZC�`�:���uX�/�E������;�A9*<��ɉ*��{�F_�]i ��D��N8X�C�j*�u&K�N���BS�ޮ4��u�fRc����n�SH��M]��U?r_
:�Vԝ��sSQEW���D�x��<  �
5�<�񃆺֎A�B��s��?W��U#8�j&���!^1�g#Q4'B�X�N,C	i5�X5@P���qɲ�Z�vڎ�Q�Y�%]ڻK���!Z����m���f]�x����+Mo*��v���@d;�4u�,<|�o|c�T\W�-7�j$KV$��Ҝ��M(���\ˡ8�R'-m�z����r�գ��5�Lby	F�3�P�u	N�2K�0J׺�I����&{���Z���L�q�پ�Ѱ�M���j�j8��J� 0�JLc0N����^���Ĝ�d&I��&<�+|L1�;�հ�Ņ㶲0��ƍ��\�4w&1��e��;�:<MKө12ˎ@a�SV���	r����%|��Оh�p꬗\���m�	:�{<�W�<:|��������v!���}\�b`]I���6�Z���(����:����$��YK%�Pd'��K��%!�&&BP��rC31cq�r#�:ܹ]V(Z*%�:)AR�W3�D��/u����]�8'�Ue%���J
�*U�������4�"0(:g�<�`�N��x����F\+��ʯ;�p���.Ύ&�)|r\s�P��ē)���Xz�-�Y
��(>&�����y�0x����(I�GRbf��!�4%8d%�љ^�㖉�k~�9>r-^Hpe,���8���֔��NGuYg!��`��e�$׭��HP�͛�Q6@s�I��K�1s�n��o9������`h8kNF�];��i4%
i���W��S3�\���wE�`��Y&�Z} Ը�pd'3�;��
r�-dt�&���X�P�]or���G��ą
^�gG�Yk�|e�!=����'Ld)���<3��2�g ��%	`�%:	�O�޵�t<��o\L�jqrHv�[z�/ �(�	����b�*5*��ݝl�C2LN�0�qr0����jKz��y�R�SUt�:�U������P���:��c]oN���0%Ji��F�Q,�P*RN�K�Bk0]Bj��&���L��!=��=�	�N�:=�}p���ae���[BQ���\CS��h�C3�C�����C�	�%��$�9	BP�f	h0�j��v�{(1����cP�%�����Jhbkϖv]�)7K��d%:$�C�`{����Uי���&Nd��db��6�~�D��&Bwf)زj���;h2�`Y	X�7�&���ЗYlãs���ij�!��A.ݢ���D]�W.�P�2M��:�'K��r^������8V={����s,� ��5������3�ZRc��9U�2I�`'QdÙ��֧zr7���ņڧC�)����$��u��31N�7��` A�s�  ��l   ����6�   �p  Դ  Eu�   � �2mM� �k@�m��,$q�H   ��Sv�\2���]�gnP.��xB1�v���TC�2�m�b[]��s�H�m�cC9n�Z������6�s�mm[$ MP
�ƺ��d�`�U��R�� �V��������J��{S�^�1���[U<�g���27J�I�N�Q�8�BN�N�#��e�K�ъ��ܭ�ȸ`3�m�e��[m�Op[�������[��4"q�H&�H���846��JV��++�u@uu�� 僂�UWX .Wm�����M4�p�uV��5���흞�Rl���5Ҫ��p�N�\�;eV�x�yn�K#�䶮�\ڬ��:�2p����m�ew-gA�Q\h�dSu�����&r5�m�H�㎶K����K�!mm�UU0�8�Y6���N��*���@h6*����I�Ŵ m�$m���Z��>��mI�M+   �m�}� :Mk�mq'ItZ[$�   M׵�mu���ڬ���Cm���͝�VŴ   	�� ��He����(-�@,6r�X��(*��- ��ŲʵSN�
�.��v�G�Oח�/�h�����5�5l,�  [mr�I5�H�����^�6ۄ�m�@m��vӺP;$����w/b�Wf��n°mV��C�g�]����c[S�4m�u m�m!4]n	�H �\  m����:X�[@�$9��m 	u�RN[@qŴ�x��ņ[r��m $8  :�75� H  �k�o�� ��<M[�ݲ�[I'�˷d�j����*U�v!����1Su VR�ͳ�$#]]c�T�=�`� m���ڸ�m�I�  �:��5@������n۳k�2��"s9:��R$0�Uں1��]�������f�!�trKiz6��Zl�Ep[:m��� �$����]m�� �l��l�N� m�Oi-�z�@mR��[U/'Y٪$m�0 ��`�i"�^�c�$-�@�!$��`�b��l�C�d�8[@h  �n��  @  ��n ��s�$3N�,۶ -�������	�-���nm[@�    �� [m׮mG  [@ ��  �hl6�  p�V��5���覨 �(U_U|W�6� �� I�I�� �:�  6�� 9�t�e���ZUBm��^Z�W5��ij���[*U -��v�i[E��[4��&�iz�$-�8b@,����g��/[KF�M��$n�,�L`-����n�k�@������$6�ͫ`����K]6�:@�8������UZ�m:)�j��
��`��
Ի,���l�` հZ����	��	f���� ��Hm�[@�m���`e�T�ەZڮ��[r�H� ��MڂA�)�Ͷp���� ���NkZ�(L͖�8�   �Im5�[RH��E���l &̣�<�p q����� �`� 7m���[m�m�-��� p  7m���   ��޴ȡ#v�n�@:j�8� m�kX��� m�Z��Ͱ$    6ͱ!�ַ�I��hp 5� m -��I�Y%�� ����k@ ���I���]0��& �t�f��8	J˱ͣU[Q����h:�I:]�`m����` �����#�d� m� �F�Ѷ��-�m۰8mm�d��݅�1���t���]iQ��4�:�l6��v ��A��[�@l��m�+'EUj�ȻJ�fv� [@6�8 m�m%�� <ڳll�8�۳��m����5���L�Z�����7�vHӬ4�[��[m�� 8�k��  �m%�mní�n Y� �Am�N��{��w��*��<��-T�U[�� h���,2ր:G 	Kh��v��;'.P�c��P�Z��� J�+�U[���\U*��=j�W̄�:��T��N8�Iz�m-�cMV�h	��I�U�PUڪ�8�*�[��m�6� 헦Mb��j�l'D�ͤFtT�+4�*�j�s5pK+U���i;���nhڪ���m�\��-��HdY$���@���R �ZI�nͷ ����EHhiiY��y���ګ`F��`,6��!�Mn-�%f��  g�da,�9�����$��{�M='FY�L��m�k�p����]�m�;Wgx�v�-ʪ�6{���<�үSI�� ��-�8�<(��H	@��R��������(��-�ݕt]�*�@U[Sq�%Z��*���@9���RAR�(n�Fu�-.a��������pY�7C�P�ڪ�W��%�k�\@V�E    ��m�k��-��khN� �g6ڗgZt�m��Ò ��n-��	8�i���M��� m�:���i��@  �m� �i�Z�I6�[v؝$k�I��M��G9m�Zp��E�#ZnͶ ��UUP�(M�
�
�|b�-�KA!6���n�8lL�k�  ��hi    m���n-�$6�-�$H-�m[@�tSI��r�� l6� 9��m�ID � �hN��G;3l>o��Z�X+�Z�U�e�.	m�   ��`6�[@ $�t �6�Vo  N�� 	 $m�-�6���H����m��b@	r��J���t�h�!��  @ݶI�m� M6 �6�m��Ke��+mm8 kZ� �R�J���.ԪpPR�(6�Au�,S��WD����Z�6�2��UR�.� m-��6�-p[F�u�u�9����I���$m&�ƲIIl��/P� Ӷ/E�}��P�^�8p8�m&À��� ېk���,L���2ãd�s�T�,��R��J��Ҫ�T���|��mɐ���U�j���*� ��M$N�l�P
l6� C����kş]ȹ��|���bv�����ä���;V�8�!q�'ɮ�l�<me�}���Y�H���yӹ�Uj�vBƅR����9#�lY QP�j��B�jSr� -� ��ځ9�� �n� [FҮ ���� p6Z�I�����	 Ύ�b�&t�@ �  ��� 8�gi��A��mo��O�4F�fsm�m�@���֤    �b� [Am8H ��8 	�� �v�      �h5�m�6� ��]6��mt ��  �^�m�`m� �M���j�T
/5V6�t       � A�$$m��K�it���[aŴkխ��6Z�[�t�m�h�	�Ͷ  � �`6��o{�� �H��m� l� 	 [��   C^���v-���H�m �6���6��A��  m��ͤ�	  6� 8 ���  ��6  M����  �ְ�e�  ��X	l�  -��  n�K@*n�V�ݒ�2�+��9j���j�]�����T�J�V�)tkZ� �m��rP-�  H 6�[X�:%RZ�V���U�ZL�[q�KҒ �d�0�m^�6ض�8  ���3����!X�R۱ �f�i0�%�-��5[Զ�:ڶ��J��AK�T��Iv��6�8    �Lm��Klu�v��0�Lm�,�i�l��1����Vvu�m�m���U�ڪ�j�����AP�ٕ�T�Hk6�UmGj�`pk[@6�^�k$��#��V�6���\��
:�b��,PQ�l��r���{=�,����<�]T�,�-�n��@�5�ֽ.�66� �UUU�@B���VV�� m�  $     x$�o �m�m��Zn���pڶ�@m�\a�mm�t 9�ņ�l�mְ   @l  m �I��� e�   �iQpp�6Z�m&�n�       vZ  w������`R5��   	�M����Wi���m�� �` m�@�[�D�6�[h
�T ��U�
U   p�[M��m�4�n�ٶ  �T�;!=R���U*�7T�Zڠ$&�^�-�-�6�8	�� H� ���H&�[R ���> ��3*�U*�UyW�vl����P �  l-�l   �  �$�~��������DU^�֗���oe!�XB�a���?���C@>�Sj��>���RGJ�b�b��M�x"��� �0 (0�@�#�tIC	�s�Ш���h 8��J�*�)�!b�{@M�a�����)܈�*��=A<EO=Q�=�j����9�A�=�[ǚC�N x�=N#�1'MA*&��� �b�H.{ؠ����>����@@2A�$K(�H40����4�H���}��@�Q�z� ��ڂ��`��0l��@v*�E$C��z@�>'`�Px�� <U�`!�sӱP��@PpQ�D���x���8L�!&��QC����� ��&���	��J�J	�`��U��!� OE 6h��\!Y�'�8�	�J'�� x��r9�A�S�A�7���y�j�У���<�T�A �8�W��QEU���_��?(��b�̒IPe���"��
�+@�R"H��̔!�(�0�!�iZE�@���ս���y�l�ݻ��`H'A�ж�RY��ۮ5��
�l�ԝVU��˩3�W���1l̛NѻRW6j��u�Z����v�[m;��I'm�F����H��ya��w%���dY�ȸ�ȶ�v�������@���UW\�T�㇮�%�b��I��+3�2!#�g�s�m�{Aƣf����zòㇳ�mְ�Ue�m�Jr��%u�d�k��Ҭ��Z�vn��u�;3���"ѝ��Mc�Tm�3�mַR�5���PPpj�6�I����iu�+�)҇���΄��+���g���pu+g9���+����s��r��W�`�;���.��ԉ��9�-��3Oe*��5ZV�`F%��5�<�l,�֪��mqR�f�cF�FZjK(%j'.�J2�56�r(�E�V���,�s���j�V0l�v�*�&�q�zN:Sp���Ujz�xh'��6����U�)<	�Ƴ�Q��U�A���I��Q���-�ag��s�D�Qۜ`�/�$]�0�����F1��N���(NL��3�h�1��KU]J�ɰ<��Hm�zB����u�KUk�7Ɖ�,�q�/i[5��5�R���C6p�+h8R�ykju
�"Z#M-դ�Ԓ�ŧ@� �j�NѰ�n;q۴��ѩ�g8��=3�T����Oxc�秚m^{d���m��ْ;u���:{z�y��X�v�ƹm:Vڭ� �Z�
�A�1=2�c;`Tڪ��jeY`�i�KX ���2��Hm=+-,�f�P]�Kq��ic��UHu� �N��Bk(ʨL���*mp@�EU]�Ҹ�x�C��jr�A������gkCU������=�:�d�����:�������V��.`.	��
]n�� iV�������I�M��bC�&��l9�E�UUQ���5�X	U㣴��R�邑݆qq��hw5�i�e]�v�m@@T K�ww������	���������@���ڮ�{���Q?�?v��v�yR�*YT�-�U�9w�"uv��gVK���-���Ʈܫ�=c]��N��ӷm��7e��v��!�̅��lv�n��8�=��rj���!�mN*�ݙx8ˎ�m�H�k�l�&КT���5�ܐ��;nM]j�d�NY��A���1u�Z��W�l�R�r�薨��n��3�  ��N�5v�ڐ��U��[�5��uT�:���{�{��a�(�.v��|�T��@�Q1��!�E C0"�Ln]Y����:��`g|�`����V޴��[m[iۥr���ٟ�*�HT�w~���0�ۋ =��qi��#���\�9��Xwצ�{q`}ݘ5�F؝���ݩ%��;��0�ۋ ����J�{w��b���Imێ��o ｸ�>����ŀwg��fכJ���̶Cm�𛛆vݶ��yܫ ^,c{���G��wW<l��\�N7LsM7|�����9��Xv{^�{q`5��l�m�N�n�`��Y*�i!�TU	�N�N��+=su����ـ慲l���RKXvn�����<��0n�,����������x��ŀy�v`��Xv{^��f�j'ww%۹l�k 淋��7v� �f��=�n,���!.mC�NwQ�{[L�lm�\mn��[v5
��p���Ӏ��g�u�밥B|���ŀs�u����Ok�9��bv�+��I.��M׀{��X}=� ����=�LV�\R�a,�-�<�����߷#�%3
8�����lI@�1(fT 	��HF��S��}�*��w���S�X�V�www-`�L��� �}z`�� s]l��-����Mݘ7w����=�n,���J�]ڑ6��ҶV�T��YI���9v�3����ZG۫q�:;���;r��;r����$��;�����9�^�7w퍱��U�C�`������9�^�7w��q`��m��wm;m]�;u�s�z`�ܬ���`��+ =��+�-1Ю�m�ـswxr������<��+�x�� �� A�@�
'�׺�\��ʼ�FRi�6ݗv�`�+ ���X;���ŀ}IRT�����NJj5Ÿ���K�V����9��.��*��r�\Zv<�q��V���pQKn�,�v���� �}z`�ܩU_q}�+ =%#�u%N��������swr�w�L���`5��=V��Ӹ�ـswq`�L����9�^��h�MW##�	�k �}z`������9��X�6Ɵ�� ;�V��;�n,��ώ���X;�� �t��V���%%\�P5*;	t.��f�� ��
@�B�t�0(Z�5�~�����EƐ5MӨX����Gd�bR%�\����V��^VO\����X�]��@��6�*������:c�l�Į������V������8�"����nׂ)خ�ŷkm�n7\�ܝ��>��e��۰\\�Uy(v������%��YB'^�0�hL�G�/:��y���F��..`�ݦza�Ã] o=\ʽ6tp3��0\L�헥�yRx<=����̮��ٌj7��k��A(�0�����f���k�Ž����c;��k��n�`}���t�h��h�;�w.���ş��g}��{ve`=@y��i�6ӫV�`}���9�=0{^�}��i͍8X��r��4�I	/n�V�k��k� �|��n�>WZ�*t�m�n�z�V�k� ;�k�;�n,�o����ڐV�wb#r޵�q��8��ط;s�����%��c������fQݞ�j�t�WwN�T�k�wc� w�׀w��X=7^ o�4�U����r��W~y����(;sa����,�o�� �f��9�0lm�����aM�m���+ �ou`��0��^��m��ݻ��v˖�%U-�`���k�;�nV {��W�Rci;c�k ��O�zl|ۿb�=ٺ��C\j!55ⳕ(��"��m\H��-�{=��]�.i^m[�ŧ�rA@;j��t�N�ݳ ;�׀o���vn�vn�{��i͍5-�E��f������#}r,Kذ�L�ڡN-`+��]��X�7^��م*�)R�ڥ�T�/r�}�� 8h�I���7leݼ_}� ����7��X�7^ o�4�U���v�[�0�L{�ŀ{�u���z����V(�F�]�˸��Q�nwn�+���ts1\&��Nz�k�v�[\��wf����=ٺ�}�������֕�m��i��n�v�VO��")��Mp�7}�Y>��|m
�*��V�5m`^ŀw|��7}��vn��@z�lR��wwܵ�*�znC �fV����U�v���)R�W�7��b��ƚ�ݲYnY�n�q`��x������o����u�]�;�^۫�6Uݭ��	7���g�:�Ç5wY�\n<�F��#L� ���7g����Lwۋ 8h�I��n؛�'wo ݞן.�I**�J�%!����>�~ŀs�u���I5[��Gi�.[�;�^���M׀n�k�9���3T,�,qX;� ����9��z{^�z��:��m��wr�v���-`��x�=� �z`��X���*�J��y:�ln�W��՚�^�7W�	���Z�<����b�7��yѨ�d�c�q��(9�����k5�c�d�@0Ί�g���V�m�+s�9�N�+���yvB����c�#�n����9�n���=7�-˛\�q�q�.�n��x��< �m��L�ܷ-#u M����3�rV���9x0���ݩ�Ný"dn����-��!4�����ܳ�e7Ι���:ݹ{�n9XX�romck���C6��O[ʹ5��k=��ֶ��?�������L����s׺�v��ʶ����J��;�nV����9��x�{o �|��M����,�v����@�Nb��q#3tc}����P��X���˹k ����{�xww�{q`M�5�n�j;ck 9�k�%}�W����ٕ�{׺�;[�4�+K�[�.�\��1;�� ���:t�ҧj�em���v纲�S������Yww]���罶���߫����\�m�S�A]�E�`�����b��"N�	:@��ui��}��~�\�{qx�ٶ��%�q�.�ig����}���{qs}��|���4E��v�^;��{w7�is���Π5E��n⻻�$�\��q}K��ٕ[�+�}���ﾪ�uIN�aN����c�z�c�n<N8:��ٺ�؀�ݝ6�S��n����&(�܊A[�K.]�w����}���}������ڡN-h�Gq˗r��}���4����d���]J+����v�ݱ�w�Ooҹ����� �'BJ��)|a�;\�H�-_<6 ��F��%o=�-�N����6p49��s�M�1��P�#�ƦY�����H��p�
iR8�x*�����c�b� ������F��-�[2i�B37E�4af�H�FQ
��:`�	⃢ ��I�PK�V']&3AJfGF����+Y���;��`=�`� ^ 9����GH��H�J��A��J-J�&J{׾��$U ���~�\R
�o�}c��Gf�oz┉C߾���JS�����);�߾��)A���{��qJR���l�?�
��.+��f*�T��w����);�߾��)J{�{���)C߾���JS� �~9��3��y�赃%�g��Rw;&�v�n�t��1�Sv��m��]k�nW�����-ԃw׽�{ݷ����߸=JR����)JP��}��R*�~߱eR
�����'�,��ۻ�k[��)J{�{���rR�Ͼ���ԥ)��p┥'~����)N���Z��-�Wwpd�2�R]����)N���R����~��ԥ)���2�R
[�&j>�b�V����pz��;�߸qJR��}��R����k�P� a(�H�S �D��>!"wt��r���W
�K_�PL�DX��Kwr򒔤��~��ԥ!>�����~��Us}�T���eRA��n܊Zc�Xgu�n}��>�y�[]��]"˱%/W{��Fmq��aoDf��Ҕ���k�R�=���pz��;�߹�)JN���=JSHߚ>$��#��R��ʤHww�=JR����┥'~����)c=8�y��K���}�$��I4�����s��)O����R����~��ԥ)����┥~����)Os��}�˶Kq۵p�^U �AK��}��U �>�^��R����~��ԥ)����)M ��^���D��.;�v\�U©R��{�qJR��>��R���{�8�I�����JS�E>�I��f�k�þ��Y�ULX{k��Ԫ(m��7V�6��2�6f�6]��Y�=.�H��P��6ۿ�=o>>���&{��R�T�n۠N��c�� ���]����	�k�.�T2o]�f�����P9�u;�V�����X0G����n8��O��-�V�YB�/7O$X��� J�/l���Z�˲��n[�9��3������[�8�ؖ}�(㭻k�$�g����=k����Ҋkδ%�����q��T۱�V�'��#^�m�v�����߸=JR�y��8�)I�����J�]~��H*�R��3Q����p���s��)O<��R����~��ԥ)�y��┥�}���)Os�Y(���Gq˻�k*�U ����b�H��<��qJR��>��R���{�*
����O��Gl�B'wx��R;�>�\R���Ͼ��ԥ)��ÊR
_n��*�T���O���\��wN���R�?y��pz��;�߸qJR�����R��y�k�R��w�g��)�ﮉ-�ݴ��{1���ۭ��":M�t���Ӄ�63���_6wLm=|���ԥ)ߞ�ÊR��{��pz��;�=�\�	rR����~��)J~����ۻd��W嬪AT��>��r3�6�%=Ͽu�)JP����=JR����8���)<���f�oZ5�u��˗.�W
�K�~�2�R[�߱=H~���߿p�t��)I��~�\*�U/h#�'�)nEww��QJP���}��R���~��)JO���=JR�~{���)I�~z_k{�j7��o9��|��)Jw�p┥'�����)K�=�|R���Ͼ��ԥ{���A�E��̶Cm�&<���7G�[�b �=�������p��7==��9��{��)JR}�}��R���߷�)J���=JR����8�)I��T��Ԗ�����H*��oוH���Ͼ��ԥ)ߞ�ÊR��}��b�H*��4��}e�6[�+$�ʤJP���}��R���~��)��D�AHy�4	Ч �O���=JR�ۿ^U �@��km��W-��yro��)N���R����~��ԥ)w�o�R�?y��pz��>Ϗu���-۷j���H*�R�w�W
�	�3�~��)JP������)N���YT��/t>�G� ݩeۊ��&��oV��4rm�tn��Nힶv�Xw��6ݫ���/GP�ڰ���.K�\*�U#�߯*�)C�}��JS�=��)JO>��W
�K�mϤiۑ]��GwyT�J|��=@4�~{�)JRy��}��R��<��p)JO~��/�f��ޣy��s\����R���~��)JO=��=H�ҝ���)JP���}��R����Y}�7k7k[����R�R��}��R��~�߳�R�>���pz���Q8�PT:�������!�qCGoa���{�ӊR��y��{�����2��ս�ԥ)ߺ��┥+�}��JS�}���)<�߾��)O����?
7:���t�r\�$0�۵�vb5��q�Ӎ��T���v�FG/]�~?��3+{(��y�)J�����JS�}���)<�߾��JR����)UHsu��߂
尸�.K�U©'~}�+JRy��}��R���߷�#�+���+�W���&��!���t�k5��R��}��pz��.����JJ�?{���R���}���);���ϋ�Yaq�v���\*�*���^U��}���)N���R����~�p�AT��~�-�WwpQ��U��}���(�'�}���R������R��߾��)JR|��_sC�wJ�kr����eH��y�g��u�;�|��fΒDx�x���k�֣�Y����:�#,�˲ݱ��&e�떙8��J�+�����:�&�'1n�C��+�n���\]x�݀p�Nncr��]ƞ�Iͦ��\����U�K-�����Z���!�;]��Od�S����;�]H��G5z��%�J;��`��m!�\]��h�i�N��AvS�7w�{����|�v��=����S�[��:v�Ǭ�]]�n]����+�7ը	��&bfX��\�e�7�s��Ӓ������)>�߾��)J]����4��}���)Os���4U��%�r�U �AK�߾�\�TQ��3����┥�~���R���~��iJO��s>���ky��Z����R���߷�)J���=JR����8�)I�����JR��O�mH�[��$�ʤH}��ԥ)߾�ÊR��}��pz��.�~��AT�W7[i�� �[�����R���~��)JO���=JR�~����)C��}��JS����f�a���U��fG�Xqճۃ`��Pݫ���nKֻ!��d�����P�N�w�{��'�����)K�=�|R���Ͼ��ԥ)���ÊR���y}��Y�[��v9x��R
����ė�*�];>!� L
���ڻ���J���pz��;��qJR�Ͻ��©R� M�w%�n�.�U ���Ͼ��ԥ)���ÊS�T��<�����)O�߿k�R��{�_n��XoQ��[�7�s�ԥ)���ÊR��y��pz��=�^��R�� C￿~��)J_�(�����V�k[��l┥'�{���)O|׿g�(}����)Jw��p┥'�����[3e�)u�����-���n{t���t��.�8Zڍ���g	���6n(�nJ�w����)�y��┥�}���)N���R����~��ԥ)w��#>��֌�y�,�kz┥�}���� �Jy���8�)I��~��)J{�{���U U����D�⼹/1W
�����8�)I�����|��#������qJR��~��R���{�s0�KqܒZ�ZʤH){���U©Q�y��┥�}���)N���R��R���j�[r�[���U �=�=�\R���Ͼ��ԥ)���ÊR��{��pz��>�5��1�_��g*W�M�8ݡ=�n=��˓�z�x5ֆӸ[W���Kn�v[��K��H*�*��}�R��{�)JR}�}��R���}��P}R{i��UvSM1�g�JS�����)>�߾��)J^���┥�}���)K�
>�}��Q�k7oz��)JO���=JR��{���)C��}��JS�����AK�|鿾%�v���wx��R
�o���)JP���}��R���~��(L �@BHL�D�IAR�$�A$��w�-J4�	,�F9BT�`�$�`����V���p�AT�=�B�K�F�v�㗾)JP���}��R���~��)JO���=JR����)JRw��f��krhC�F����v67m;uI�S^�WSЅg�q�iR���;��_6�+m=|���ԥ)���ÊR��}��pz��=�=�\�2������ԥ)���30r�w$�����R
^�~�p_��$2S����┥�����ԥ)���,�AT��|�}i�v�,�.X��=JR����)JP���}��C�f����ÊR������R���D��n�v[��K��H*�*�}�ث���{�)JRy��}��R��J��y�r��q�6
��4�I]�w���)Jw��p┥'^}���)Os�~��(|��~��)Jh������(�%���#)�M@�/B`0�*i�/4a��U�8d.E�#��L0���C)CZS2@E$,QHPĥ%A$��}�f���1jg<l��$$�	%kV��6S�JUѶ$�`�����D"tt+�LR�:4卐rx�Be��tc`J��1'f��"�m �ZR��)���("s�$ejZ�$�������&Id��1��5��)	�A�m��
��N�!K5�	,!!Vx�b�}��� �Z�a)�M����Z]5h��0�8#4q|��uK,O<N	!$AT�Cp��ݝ�GP��<Ў&�c(�D��
�8Đ���L��w����I��� ��f$��J�Cx��'h�I	!f	R�	d
Ifd$ �a�Б���.���z��VY��[�;��A6b� b�fD�-��]EhSC
�+22�B��L��M2l�t$R�/ƾ��֭tk7�ᆳ4u�G�5���J�jP�(��4� �m��,�f�@;�ߵx��ѳ#�7�m���8@�X���뜩�����7M�-��Ϸ<WG;XM�� �#������&;>z���-�&�n��[cT��&����w[˛n7<O�h�$12Y�3�q;�ۍ��f�ݞ���ð��nWl�C��ݖ�q��R��3�\4�0ݖ�g��.��������Mјy^��*����]���*F��R��F���մ��:C���&Z�7eX
U]��SOe��c�+���5�M���{\��T!�Ð}�z�ٗ�j�x��^��Y5��0��ևF��� �)jS4�$s��Tn��SQ����+eRT:j�+B%'d)0CRJ�Ԁ��@�J�����9B�TB`����v��vj�r��=��$��L��b�h�h-Б5��P�H�b����|����P��I��������Hk{Rd&�v��du�كO=&D��WS��V��+Xv�#R��
z�A���;`�{/k(�gnc1�ٚN�pu@:������U[��������B��K�*����T���%�X[ӟVi8�����z4@r&�!�b�;&�^VԤJ���:!�q�meN����eȹx*����x�#��C����+�CG\غ�6��x�kג�ĺ�`+���L���	�����X�k[f���BR:i�*��xȬ�̩W��^5bI�i�h�*��� E�Fj��ƪ�� ���Kv ��_��핛E�T-��U�UGa6��iV��t�*�N�lYv�u� �bh+� U�2�ɻ7l1/k	N�y��2��b{y��_Y6趂(�L�z���휾�ԓ']=im]S�ۋ��^����sj�;A��h
�j�Wv�^ݻj�̲#��m�]5 ��f���$'�\v�JK*o�.��~+(*�T��1��ß*�D
��c���}����N�נ��סاh?�ôPN�1��('�6�e�{��k5��Z�"�����n5p`a�v��rp�T�����b,�U�Ya��)p���f��F�����R�^��x8�u�A�ω7�_mds�[���S�i����ґ�q���Vs4�f6��"��V�=�xҸ��7Z�WT��Р�)�����Ƽ�;d�r��vB�y2r[��l�)�c*��U�Ʒ�8W�m�tE��=�۰�[���}��q@�kv����BW���ܼ��^v�{#Ӷ�b�v�1�Z{�ܡ;nԈ�mp�Ieܵ��R
^����ԥ)�y��┥�����)k�fV}��P}S��)t�T��Qm�R��������~���R���߸qJR�����R�����5������.�R[�߱W%)N���R���d������)��cy�9�r9�P�n�"�����Z����R���߸qJR�����R����k�R�>��pz��=���d�;j�ڻ���R
\���*�)�y��┥�����)N���YT��-�G�(�����-��;\j
=��6�Fd�2�)�S�[%�nCq�\6�.K��W
�K_��H*�*��fW�*�;6e`����(�q'ue�-��%��5��}|�)i��X�MRF�I %�t�z �κ�����݁���Ȅ���UM(�4��<|ߧ���9�5{e��� �������V�v� ���X��z/��Xo#�^׷}�ݔ�mRC��m�j���
�;�>ٳ+ �ݜ���wJ����,lD��n&7 �v;BJ7 v�������9ȇ����mQYv�ҡ�ջ�"���f��@��;�DG �����sP��PX��;�yw��f̬��vs�j���5wv>~H�Ti
��Wwv�`��@�[۰1{��=\�\�Y޺�>y2���4�v�v�5o��T���x^����2�;B�٘w�ĜP��wp	w0>�f�R����9���W�^��v���)�M�*���p0���a�U#��c{Y5�vtv��w7n��aMS�Ht7mU��I�<�|�fVɻ9�5{e��� ������M���e�u�s�g8�l�˻��͙Y@OC䤴�А�*�|����.���͏ ��p��EK�uv�A
���5d��� ����~x��y@|�2��H?���nш�j��z�5j	P1Sٚ��fǀs�g8�l���l�&�n}���L��ku���n�n��mڹ�\.�p��v�㱺��k��^waa9U*��x;�s�j���;��ˮ vlx�x$t��V;�hv��;��`��e��������(�q'vU�4ݖ�k ��/�ݏ ��9�;��`S�H�[�uj���O�2�������k�ޟc�=8�J��QS2M%5U�/�n���:z�d��uUߞ��U�"���`��N�Fb���{��]��=��q��K�%l��͑��[\��I!����
�m6e�zuls�Ѫ ����c)�R�ѳ&��9�S��r�yzȍ&'*
�綧�Gb\�Ȧ���N��	w�WC�u�#��)Zi#7��u���yՋ�;����FŧS��<n�AԹ��@Β��F�R�ZX���m�Ի/J�Uw�F�r޴����RM� ��%��$�e/Nq2��Mr�r+���%����pXv��z�쵺�ۈ�q�كi�����R�
�$*�UU~~�k�{'� �1��D\ ��۰��512�R�qT�������c��{�vޖ�@9�BDQ���W�������n��-���nl̔��2L��iۻo ��9�;�`��/�Q�lx�x$`�۰�ݻ��� �E�?k�/��ݒs�z��U�����M�{�nx7=��^�M��֣��ք����狞��+۫|�w%���6����/��ǀwd���Ȱ��T��r]�,�^d���ד��Ui(�MՍ݁�Kk�}��9��r"@NƩSU3$ҩ������������e�ޑ�!�[,t6��aj�������=��̀{��CW���`=PF����QJ��SK�{'� ��xvI��\� ��m���T�ݶ��xӱ;n��X�=��7X,��ڍ���67m���)f&Б�i&��O���c�>����mtd�s`>d�&虒eL�*����cn�y�9Ȅ�9�]=9���۱��(���Ac�wM7�ݹ�ߤ��nͽ� �������Օi�7ai��{��/�� ���7��OW@q���4�dUU7l9o/�� �f�p�ذv�$��*^����	"?�%�m�-��\�6�R��nC˵�X7�aӵ�\���V	�$T�*B���׷`|���|��}���|��:-���|���`��K��c�9ٳ� ����n��*i���ݿl� o�<��9�;/b�z!"KH����;˷�a��s��ǵ�>�{v�q�����9�R����UUs��������~��ԒI-;�m���s�uM��qwv> o�<y������&��STQP�swS�]GB��u'4n�n;66��&;��j�Z݅�[�+}�_���8�� 7��{g8�Q[W��Li��ۼ����}����s��*{i�V[���q7����������r8��{=�����'$I3I�[x�s�E헀qI��{c�9�>JK�HwB��8^�xx����@��;�/�|#����gƞ����<ڜth��t�����u�,s�==q�N��4km�̛��\�+��Dp@Dx�	������EٌuT��.�p�&�[n����MМ�����y��h����%:ݔn��FڭH�m^NV�v�'\*��m)ՠ
ӝ�iG2E�SJ�7V{Ncq��&U,�eҽ�f���ø�^ѐ�l֒F6��kn�S��a�nu��`h:g��gs�mu�Og`�#[!nݶ��\,^���S9w�v2ćDoL����j���@��;��9�.�!#e�X�`��]�> Olx�݀ױ�@��:��$l9H�UR�I�6�i6�&���^�x� ;��T�c�V��Xݻ�8��^i�u`y��lq7�~�=�ⴥ%ZcM�bn�M�8�H�	6Np��]y��pL�"TLl�3RUH�}�z�Sv���]v�n���� s��w	�q��iYnӫ}M�g@=��<M�� ��< �d�����!����xx��"}�Q��9���}��7���� �ڤ�X�m	�V�� =� $�3�P� �d� =�"�m;J�h�]��l���G�OI9�*�{c�:��	-"�cVb����c�
�zI���/ �vGͷ����}��!�zz�UoM�ǓX�;���ڀ�jCOY�~׾O�;<gw�����9J�T�*������`|��zY���r*��l����O�Ҷ���mݴ�8W�^쏀� ��s��Em\Yi�7v�w�E�#�}#���>�[�E�I�qT�"����6�hrF��Sa&n]@�Jv�PF��D0ΰ�`v$�z*��qU��D�dI�	�I�JQR'��ػh�h!��5�ֈR�MtXF�7��LNל��>;v��:R4 �� w� �@zP4���Q�D�b l��A��i�s�@N�=���b/H
�;����Uy����W��R*1���i�g�| �x�'8�{�>���JXҫ�wt�Wm�I9�=�ذ��������R�����.�Z�����
r�-����>{�\�6�˜���݁vg	��/p2]�E$;m��n����H��H�	�Np�R*vӱ4|���E�G��G�M�s�{ױ`]�Ѝ�*���U��c�}#�&�9��|��]S�ڰd�9sJjE*j�)*��	$����XRH��K�����j�v;�v;|���XR7V�����n�|�Gf%)��3��z�96�ݡ��s�cƛA�m�x5ъ�p/[U��HD14L�E)��U+ �{���G�I�s��^ŀz�ґQ�aWm'c\o1����	6Np��,)�>���N���wt�V��$�9�;�ذ��| �<݊�R$�t$;�v�� ���,)� ;� ��s���m;�G��XO1Ձ���v��n݁�N5�=�� �@�qZ�G�&8hE��L�ɈH���K�Q�:f)	T��A�`�E1�s X���paH����NF��k���Yx�0���pp�[&uv��kj�Ԯ��/�n�Qg�JI���e��A�{S�ψ��9H�`��n.�)�(m���O=gP�6�Qcab��8؊���d��d�v�n�r�dk˻=��1��^Ņ��Ѣ�
!=�H��(c/)tu����2�5����z}���|��X��87g��2;N�SL[���3�Oﻻ�����ˡu����nu��Yݡ�X�i�8�{@<�nc���dƾ8�N�"N��k����~n�zq����u�%m�K��ݗj�i��x�����>z�,)� ;�G������T"J�UU]��k��>����G����v��A-)*)MI)6��vg ;���9�+޽� ڞ�D�:���C\������ս�3�{ױ`Sv>٩L��Ϙ��3^7� ��l:x�s�[�b�v���o[ϞͶ�"	v�%�)m�w�ow��=�ذ���\ �x�TW-7m�#e��{�~x֤���K�T�$�v"<�[�`u�@ϱ����p�T��4��v��7c�}��ݓ���� �[Uc���1c���%�������¨��{_ ���m���.�ݱ�m�{�s�{ױ`f�� w�<IF��N��/w^�r��l���Ƈ��J<�c.%�v�V�\8��N{_*-ݺ�tݼ���Xٻ3��ǀovNpx��ږRIScBJ���ٜ �<{�s�wױg�mvm)���Wm���p���ݓ�5����%�\ \!RBT2E;��W����Uu������%)4��j��N��7�'8�{ vn��Q�H�v*��Zn�¦�!���헀Wf�� w�<{�s�w��$]T���j��+t���Vg��ᗷ0���p��7<p��˟#���r�vZ)���ۼ �ݙ��G�ovK��1c����D'�)(�
'�v�� �<{�s�u{e�f��+m*�jحZ�;M��ovNp���(;7fp������+m�"�N�j�7�
2q������>�u�Ȉ��{~�pz��|��ܸ(�� ;7fp
;���9�<���֒L���4p�b��s6;pv�ڡ�:A/ӥ%�gC��X�T���Fr�L�+%�Z�ݼ�5���n�}�݁��s�h<��������&jT��UU]>���p�c�:��| �<���b����(@��6���c�:��| �<{�s���*�S��M4S.�����n���c�7�'8UQ�lx�t�T�����VbǏ��ǀ~���w�y���\����~�UqD܈�����������o#�ⱚ3�vu�[]`��6m�WLkE�#�M�b�n�۵ìe�ה��v�<<����iv�-��� l��U�71�]��vPv�c���Q�V�fE�9�Q�m�Z�ݺ���.�:�2�S��Ss���'dJ�RKqQLj<V'ێNԧ��n�x`�Qe7�D�|ӵ �fsez1Y.��!	�
z��G*�8�����ؙo�����ww|�F�ۏ����z�IH����n{{m��-�l�v��; &X�Z-RM�T'�d�H�[�m����8W�^�7c�}��^�7n��wcV��:����9� �������}�ݜ��@w��&��&5n�w�uM���lx�d� ����6�6���ucce��o �����������헁�8DDqyk{V�	5	*�UIU7�ovNp�l� �ݙ��G�{�����m/N1n%��oomlt�m��[,��uN\���+��,����v/w���f�!����/ ;7fp���直��� zK���N�E4��w���9�?"1��^���ʺ�߾못�=�\�.�h������W�c��}���7vj^X�z���`8�Jܓ,�V��Ӷ�>�����^�xTݏ�}U��lx��E	�wH�Ӻn�����@�Dzu���=�k�g���Kw�"�iݻ".\M0����nۣui|	q�$�8s�;�h�z3�>w���j�����[����Sv> w���9�:����͠��[�:���cx��ly_}@ovNp�l��n�����R���um&��9�'8W�^��RDL�+����{�> {dx�TQ66�J��-��Ȉ�{��f:��������~���6uRJQ�������y�����c�7�'8W�^=~ۧ��e�eXA�]t��\�۷cp�n	ɱ`�)q��n��18bJ�db���wc������lx�d� ����:��|V�T),�eڻm4���ovNs�UR��Z�z���`{tf	�
�jam�7o���/ ꛱����c�7�'8}@l�N�ZLi�V&��n�����߷ʽ�߾��S���#E
/A 8p>=AG��}�r�N�PJv����cx��lx�UP��{�X�z��:�>MA�DȢY[gbᗛ�㣊G�ې��v{@r���|�+��	�������x�I��헀yM����}���UF�lv�J���m�u{e����7c�}������G! �\#gU$�*��3S�16���c��s�^6���{��ah��J�bt]Y�3�UU%ퟞ�׷`|��zȃ�=����	�l�V��I�x6l� ����<��7�W~{��W���i=�nϸL�?ǘ��AH�)�Rվ k�+�q8��Ju��3��W:3|SÛ��F��@l��0���~Aء��}�"HH� � ����"Z	"!��@�^�r3���9��������٩��a��;()(a�b�ܻ��Dwl�Xs��1"����Zj����`�B� >&�F�ɉK�f-�1*q�ą6	*��5�
ldٚS� $%_�6Y� v�B�i;�HP�%"V����b^�:�3��I'��v��FK�R�ր���z�Ŗ�m�"��׫2l�EۖO�i&kɸf���-�bv,)Z-Cĸ��Z�h�i��\ۛ!����;��g�½n;tȾ�t�V�ǇER�����Vʫ e�vrm�� ����`���h9 ���v�&�/�]w�ltv�"5��7U��G��]v��ŲD��=;[*���Mv���R��k�Mpa�n�u��[=6�v��<�Upp��[x�U�WXv�� v�t]��݄6�L�t�.{\m�MM[U: ���(pY�;������&�`s�\���.���i�O+�W��P��:�v�ƃ�t�rKw:���\��ɳȚn�V�2bp�691u.4�$h*(���U�m�&Z��J�p��*�q��,�*�$&�
�mb����*�\4H&�J�G2�<8�QT<NL�-�;m]�;�<�$��"L���E�Aԅ�e�!��S��L�+&֛���瓪�u)��K������tsj�q����\JЬ����1:���vw4�R����[��U��%��q�A�ŷ[[����OH���og��A5Y�:ve�- �Vܰ�+m�+�wi�w�;sFY%o6� �GSJ�URe�V	w9�qa6��%6�Ry���e[zN	�G8�5&��^R�n����d�y�2M�l;��%�5�$)\������3ف��8�u���Z����͗v:���u�y:�M�ڤ��u<�vznX%�*�j�J��ky�X�g(A�s�B�0g $ؒ��T��Ey��u7@�I*��y�4�6������k-�mZ�m�֛�m��I�E[��eEژ��2nSyǭ�m��b�n�� ��2� ˳D�W�`g���v��!��F'��v�Wj%;v;<��:��-�u���І�
�UV0��[GUK6F؃�k��\ *%"]�٩��J�Mm��:*���+n8b�B�V�$�H�@�y�vu� R�5w����}�ǫ�����}��y�!�t(�����h�x	�}��ا��FtkF�,��(�U-��=��9`1�r;`�֛�2�Kz76M�<��'�Q��A�;�;l�et�n�9�o>:��A�9fӄ���Ҏ�m��`q�������:��Ʒw\�l��Vp����v�M�[�V�hS�F`�sۃV�g��^��um�ժܘ�]��"�<��y8�vԝ�AZ�ٔ3�PVE�Q^I�VI�e��쎞{��v�Ӿn�Řt7ZH67Dn������͋����)N�v@��pX�J�ݻ�;n�nt�K�<�� ;� �͜��̧wV�ƛ�bn�)폀�ǀof�p�l�k�PJeۦ[-�cx��H�����^ŀyOl|}Ap*ƕ�N���x�l� �b�<��> w�<�ʩl���¢��� ���O1Հ}��gͻ�6#���o�u�\��-'L=�l�tm�8�t���WK��BIyC��ݕ�8��=�b5��*iX��� ���@ϛw��|�2^������V�N�t�1����~�p�C;��r9�"���v�8�@�y��b#��P(݉TL��)RUU]绷`{Ӎt,�u`y���bN�j������8�럖�I�����l����5��դ1�vZM��wc��U���쓜��� �|��D�
5>�Ip�B]�-�e�$���]]�n]�繶t�SI�M9�W��L�!�_j�V���@�m݁���G.bm�X 6�KbJJ�IUUt�����X�����c��ʩl�������8}7�y���Ô�T�K8s�苻'��|�<P�e�$�TʅSK���oj�=�k�^6��;�ذ��K%
����f> w�͒s�wױ`[� 쭙�5�3�k:��H�>k=������n��������㓾?;v8�c&�7E�[�
��绷`}�ƺ�f:��������J������8}{廮��c��xۻ��${ :�B�����@��ڰ���o9��%��۰=�?,Wd����1ն�\����c��x�݁���"#W!p�,!��@x���,Ͻ������{�K�X�eӫi6�͛9�;�ذ-�:�����s�����TT(�����wV��d�;��o�֌�,�Ol��֍ܛ%���.�O-]�X���y�=��� ��l| �<�6s�-)Uܦ��LrH�it,�:���r"!s������g�p��,��B��m�Į�fU�}�u�/;���}�ƺ�{XKT��jح+t���6s�wױ`[폀UU�ǀI��JWn�cwm[|���X��c�}��ٿs�]W�T��R�J�>�Y-�8Ki��6^*Nݺ���� ī���a�F���%X�Ru�&��Ŭ�s�4�c������ӱmO5�21����B�Q���m���9�k�����#��-ѽQ��a���gQnD��[7'"dx	 r����q��[���NW�m��2� M��!>[�9�ڱQ��cY��JQA�[s�{*�U�C�4n�)���%�(�\�KRꤪB�JS���v\���vh��w�;lc4v76���3M�ζ�6���e���wo ������]��9�>�/W@����$��*&isڮ��>�:��9��׷`{%�����g"9��rE%Dëi6�͛9�:�����$o�< ���=�ilRSM��`	U$��� ���������^݀6��.)9�I���߯�*J����9�g8}{��IJ�vU؝�X�.�>nn:��k���z5��k�㮝ڮU�]���ɓ��V�t���}��ٳ���kb#��DD Ÿ��d��j�j�)KW-��x7���⤗˕J�R���>���7V���t�r!���UA ����p-�� ���bG}�����8|��j|�e�v�.�R_S� ;� �͜�^�x�IA��KVI�|�/3���x~o�uI/l���g��c��ğfk�P��:�5�pX�o.;x��#��NK��ۙ�nv�6�"�XҲ�մ�o ��9�:���ۻ3��H�l۪Q�bo�P)�5W`{'��ă5��q#�v��|�v��∄�H[T��jR�T�޷�����Ϊ���˰<��v���j��۞�8v�,���II[ci)��v�����t����ƺ�,��Ձ�JKv���*Jj*i*���xۻ9�k�yfc� ���ۃ8�0?|�Չs��M�L���1��ƌs��ˉ����\v�ll��[vթao���ذ-ݏ�ݏ(l����2*%�e*)R�5SG@���W��q �{]绷`}�L��|��D�EJ��m;�<��I���'8w\0-ݏ�{��}jƕ�N���x6I�U߾��^{�s��y(���.�����m�(��o�,�o����fc�}��^6���#2AHq�
��7|g���,�g�ZAӚ���f7`��֠}��uRK*�����m���_���wc�9�NUp��xa~�.�(Vݲ�щffp����'8V잁噎�c���.G"�J[�UR*�T�U5]绷`|��؈��6���?<MJRN�����Wo������s�<�1Հ}�u��G"!|�w�� qQ;ɔ��UMT�,�u`o �r8���@����,�=!��A�&o�ϖF��G�[^K����=\��<���ƭ��t�6L��jzxX*{#8���vy�0u�e�=����v�FI5(h8�;
�5o`��.�n.ի>�9�Z���ֶ��4&.fH잎�!vQ��D1�ܷ���Vvɮ�}�u�콵�u�;�s�=��.v[.���x�B��kd�YS���D��:;f��s��N�U0�3f�e�n�o[�{�A������}o�����q!5Ь���<w�j�mW;[W�x1�,=�۳{p���V�n�,i���| ���sd��[��ꪠ<�v>���3�V4��um+m��'8���-ݏ�ݏ+婢�ͺ�)*�)�$��� �1�@���V�8��Ձ��۰x�uU*�jff)J�3U�<�v> wv<�$� ��㻱����%JV��j�1fc�wc�9�Np���[� ٴ�]RU���f����蹕�r`�ݻm���`x�\���8�Ǭ]v�vm^}TXг-ݻ�i6;i&�͒s�f:�Y��y <��@�`����]�r[�����y䫂JĄ�P 
z��`�~�t����u`cu�/wz�� 8���Ți���j�~| ��xQ͛9��ǀwv�@��N�vݫ\ǘ���]�� �1�Cc�'�j�y�����J*&�������^o_ �6~| ��x����VZV]J�oNtC���n�q�}۔�S	u�Fֵ��;i-�Eoc{��3"F]���I������=������l�� CuT���v��ݦ���<�����x6l� ;��_�����ڶ�1fc�wc����~��<QD�R�4����QE1�}w���&3a�l�i)�I�£��޺�oB�����u��sm�zs��$�#.htFU�pu���\�����PD���vP;L5.���M�܆I���p�eA�������hf����LX�A3О���F��\�:⚚ ��F��P:h���sG��X=
T�Q,#�s�����{���P�F/ IR�
�T�� zj��( �0ثꨤ���A��'���FOajj���-���&��%��wm&�m%U]�s�!|���M��,�:��c�&�+�鲐�ݱ[� �ݗ�69�\������tǎ���q/|��Cx�;v�,�[x	v�V�n�Bs��Q{l����DC�~������l�Ͼ�[����Hv��.�j�� ;�͛9�:�e���3���	N�jƕ�[J�x6l� ;� {}�8���mz]QM�j�]�� �;� y��Ϊ��߷���>�1$:U;�����=.{xءR�cM���V��o =�ٜ ��x6l� �ݗ�~���w�����׿
�B�[��c�]d5�n��Ds`C)S@�tZv�p�%v;���N\M�N�K33����9�g8V� ��fp	�����j؛��o �͜�_Pun��o�g ;�6@�]'M��ƛJ�8v�,V�c���@wv<�l� ��N�}v&�i��T��DBr��X����;�#��}��`ݠ�E]�v�����y���u�7��G>�{��y���1g�Ձ��w}~w�����Ɔ����qS���7>�gD�\p��_��\��������ȶΎ�J�A�]���A���;]�㔩���@�!�
�wWK,�\�2:�K��M�k[�x�n�,�#��m�M]����ƴ����Kc���;i��Zy݆�uEы.v�:�앴�m#V��\�2���[�T��I��y��y}����)y	t��=�����~{�ߜ��^���}'��h�����}u�p�^�z��յ�$��]�����"����*R�b�yV�Wt�[I��	��9�5{e��� ;6<ҽ.���&��B.��j�9����b9 =�k�}���b"#�9ȈA�2������U!T�O@i�ڰ�:�}������5}�d�:��5*h*�GW{ڰ9�������^�x����7KQYwe�6;i+o �9�*���V�V�c�d� �J�
�N�e�[e&�_Ȩ�X��ͪ�..t[q�wD��;nݓtt������]sZ�����|��e�o�> vlx���ݠ6�FUؚhlE�x[�o�;#昅�vzN�]WǀMݜ����͠�*���vݫ|o1��c�'f�p���5{e�o�>=A)��[]�um&����{^�`5�g�5��V9�>x�yǜ����֨V��8�l�-���͏ ��9��������B�n�;i��g:��9���G�m���q��8�r`A�:n�n�[���w�E���ٱ����E����^�Z&���V,�| ���I��W�^�}�����-�ڻV��i+o �9�5{e��믋5nl| �����ʴ�I���I�p�W�^�}���c�9&�p�өL�M��� վ��ٱ��g8�l��ԕR[�4��$B�E��c�p���NƷc��t���v쉷n�j�F���o��z����Ԍlm����@=�~x�����/ �}��	��b�մ�o �<wds����5��V��]��G3c\�-�)*�J�����ǳ��c�W�fǀN͜�ե��۲��;�xR�� ;6<vl�~��}�A�T���-~���_{_�P"-��4�Y��ٱ��}�N͙�5{e�o�>��-�V]';���z�xy�L�6�'��l��v�l~�;�;w���۴R��ID���RUM$����k۰1{�����#�Dr9���t�[Am�m4�ƛ� �헀E���ٿ^�~߹�I~J%U���Q)�A9%��ڰ�&���e����@lN�N����-�> vH�	ٳ� ���*�"�l|z����N�N���vl� 7v<-���� �UI-�V��(�"�M�bwa-7wb])@�Jv�/렇��i{Y�Y�����:&c]Q{=8�ݜ�v��2�v��[���u�R���b���<��P��z-�aa�:�ډ�Ҳ�Zv�H�l�#�h2α[~t	�At��u�g�
l�m]ª�t.�hg��#��¤��t�vd�l���0����ZF��Gx��[���]��f���c��{D��{���?Wϩ�mu�JuR���x��t��x��Y3زq=��S�M�\�=���#�z�66�j�e�� o�<-���͏ ��9�	�J%7V�E]�����o�> vlx��� o�<�EU �,ۤ��Lm�N�ř���?<vc�5!����=�0�!â��*iT�J����[�{vX�zY�o���CR�E�U��o�W�^�c�fǀN͜�,Y�P�枞ʛF�L�[o8tq�v68�u���lsb�5b��XSyJ�e�V;�K.�[w�E���ٱ��g8���͠��'L��mݾ[�| ��}�k�����k�� I#�"�l|z��IB�ub�V�m�vl� 7������X��t|�� uQU\�	E5vȈ��9�=����ڰ�:��g85V�)�v�v��ۼ-�:�69�p�s�^׵�7���=������s�AH[˴�v(�hb���Y�ѡ��s�D�w�����P/;��������:U�> vlx�����/ �}����-(Ʈ�V��I6�	ٳ�*��}��o�> vlx�IjW(�2Չ�7� o�<-����WJ t��� �`M{;eЫ C2�%@ĕ��C���ҀHA!*�o?)򾂉��~����9�7�:���E���m���^=� �����x����s�>y l�-���o�� ;6<�W�WԢ"""7��� �=���{X�ى��]��[��hޱ���q�5Q�$tX6������a���v�u�_X���^�=��:���9��]ݔ��#t���J�v��5{e�"�c� �㮀�x���Ȅ�Z�N�PT�,i�ۼ�?> vH�+ꪪ�vl� ջ/ �#�Ii��n�tV,x��#�'f�p[��=�R���}�ETWT�Q�߯�wco���[�ۻ����N͜��e�o�> vH���
���V�I�YL���SM�Tu��pq�V���r8q6��n���ÎK @ܭ�I��7��v^�c�d�>���	ٳ��@h�1��H�� �}���G�N͜��e�W�P�@lӴ��N��| ���g8��x[폀OP\)(P��N��櫡�[�{���{=��:��.G!{wk�g����ffyJ�5v,�=��:��������>GB�r'9H�R�����CF���ݤ�@�])�C��'��l��A<���b0�0dƔK�u�[S�b��R�P�П!9�Mf�ȱk�D��CKEMD�����fZ�Y����IJǆ�4+Ლ
Գ�t�dd�����b�"
��(J�p����� )%��,T234���-5BP���=S�r)(B00��JAx�x�fI2VK�g@��pA�T�Q&�%T�c�B㻷q��ݷd���N�����umm[I��\�`W�r��`'\�3�Mr۲�m��W]�I�͚�tFJ
��Bkh������Z��qdm�a.s��p�>-��n��d�5V���T�s��4Fv\�]X���x_V�/R8r��-u;r�R4��m
y��Vݛ����c�F��v۲d5�N�j���Z��)�۵�=z��qPm��T���r@�#M�vѳ�p ��EӠ�,8�e٣�9[�� i���4]ZgW�$GT�1��6���C�-)��c]zm>T��O�P5�]@x̓���ݢaݻl�vN+m��"U[fqIN��Ms�Z�9}�ڣn�'b�nP��U�.T*mF�eSzWD�U���D�Um��@ɒ
U.%D��ٵb���F�)��D�c�R�v^wh^�"��U�q��j;v7k�@5U�]�e�^M�Egd쉍��S�gz5ȼ����X��E�ۚ2��T�����j�S�*�-+B�O�6n;L�'S0��M�����j}���M��=;֏Ii�Q�k����W�F�:n-Wl�Yi�
��4�b�̅'d@��^��;4��%aԛA�΃�@ꪓ'��I�W'@�mcuU��R��Pl\�5�71����`��lxt�\�-���%皭��\�ɪz7K�5Gd=��SK%��$غKz�9���=���&�qQ���v�.w%�ؚݸ���K��燠�P�u2��/m�i�qY�]Xʭ.w%mtm�m X 2��kQ�ܐ��뽴���V�A�d�	-tki{NiZ�鶕UjR[m�$���m�!�Jt�Aj�����V��S<j����s�rET���4.�: We�ـj���u�ή��`��L���zT5M�����Y6.��ceN ��x*�Z�� �.�[+% /EZ�k���SW:bk3 R��n�+��R��[ T�9,��rm[T��x;g#u�ځ7n6�s:U�����{��t��F��{��*�����hb��x�Ҟi](	mRT�����WR����n\��v�w:����n��6�G�7c%ͼt�]ęy��J\OZ݆ݍR�V<f��挽�Y��i�sϒ�dL�/2��{)�&�����:���Y�.m�]��� ���#�c��9�9��+�7X5��i��b˵����������\Ų9�ї����vn
�
�S�z��Mϳ��ӌq�n7Y���j�v�u�C3�6|�-���]��ʆ��F�#qh9�v��ŕNs�dA���93ؒ֬�x-U��cM�cui;�p.� ;�W@<w��8DD|&�z|��	��M���X���vG�N͜�[�����Ԓ���j���v�;6s�yn��"�l| ������:%TQE)���c������@���X��t"��vd(�RT�cb-��"�l| ���	ٳ��v^��IV��N���Qm�
�J�m�q��E�ţn6�v5��>����m���m���m7n��| ���	ٳ� ���9h5<{V��	i�ED�J������J����U*�,n�x_w~� wdy@{��Ļ���K�E�� =��c�vG�N͜��Jm�7e�էwm�o�> wdx���G�c�8����)&�N��]bǎ�>��lr#��׿|��t���Ϳ;�ߟ��>6G�;%�*�E��.�=v;o=�m�άJ<Ҧ�؛]�ۜ]v�v�\ u$�J��i*��}�n�=��5��Vݑ�u*��鍥e����nǀE���ݑ��Np�T��h��v�+m�n�| ���ﶢ� �P� �Q)De$��Ab�%q��9�{�g8=#�96���m7n��vȀ����m݀{1�Cb���`n@N���Q*TM$���?�w`ݏ �wc�vG�{����bJ˨�:p�ɏ]cr`�g�s��F��CoI�/�3�����L�E�%[Mբ]������:����Dr�o�v�qF�TR����ӻ���v> wdx쓜 ��xWVд"i۱�V,x��n���vo1������`fJI	ԧwm'M�I�x쓜 ��x[�PUW>�UW�WLS#�9tD���i��cV��nǀE����#�'d�������(��&6����|�lݶ��t�9���-ۈ��kL��;l��M��V��"���ݑ��NW =�ɴ�Ս�ݷ|o1��n������݀c{]��u{
�:BZRB����Ut��݀{����s����Հ{7k�{�	���fyJ�A5Wa��q,ǵ�56���7]��D����L!�Δ��Q*���5]��:�6"#����`o�v��=�|�`��GX(��Bo-���닭��HJbqs<�Vˎ�c��<�m͵g���"�O&��Y��Z+��(8^�"��^8	��5n�=n����&�\�r�/N���Ok�c#�X����Mn�f��v{t�c�8s�C����ڨ�"��9<l��a��|����q�{vz�6�7U��[`k\M�D�s�k�^S��H�^Ґ��s<N4*�8��I{Ivƚi�w��ݽ����^������s]��l+�����h���N8Ƈy�;���?����tT�Tuv�L?6��� �c��g�>�i%�۴�lvһo ��9�nǀE���ݑ�t�(t��e�nӷ� {v<W�#��ݑ�������i4P[i�V��5{���${��=��v#��t� �մ۷m��| ����I� {1�@��7VǤ��\S
'JEL�rbn�ct��,�h��b��七c��������
�)J�I*��=��v�c�W�#���ݑ���K�e5Iձ�� ���gˉR�I*^j���~� zlx}6s�<�n�vեi�Iݻ�<��> wdx�|w�g8��T[Km(�lun�
�� ;�<��9�<�e�]� ݴ�JF�I�cv�v��M��_U}�/ ����ݑ���WwR�j����(���^�˻ O[���t�jh�v�����;��Rt[��e�n�[� �ݗ�u{d| ����d� ��i2��Qi�iU=��n�c��DB��r9<�k�{�p-�x��Q�մ۷m��|*�߾�*�Ͼ���� �I��8�Q������ֹWY�߾�U}�__��jԶ���UU*�G}��8�ߞ����#�=�J%�j�`�Wv��nǀq{d| ����vs������:�]v����[��R!���:uV�zNN�;r����x�Uy���w{���I�>Q���+MZwv�����#�;��� {v<T[JZ��m:t�.�<���%}U_W�=�f {v< �^~�Hݴ�$n��i�ݴ���{d�� {v<��#�vG�mMҔ�v&�
I��Uv�Ȉ�,ok�|��Հ}��A��@r=�9X���`�n�nڥm��}#�vG�w}��َ��"""9�j�&f�!4�����],3���۰�7[�Bݹ�V�X9�C뺓���%� 1L�r��˗s.�/��v���w`�u�-g�����@�N�$��7�'8����� ;�<�����=�J%�j�t�CI�� =��7c�vG�ovNp*F�ݵj��C����� ;�<{�s�}_UWǷc�<����-+lt�۫�O1��#�7�'8����߯�z�*�"5��⍎���A����� /F�9x�J[���sI�����t�4������2���݀��ѣh�v�s��(
���"y�MN�')�*�ԇ#��O5n�5ۇ��q�"��˫�;#(/i��/b��Y=�o�vCv6����n�}y�[J����[O:8A.�j�`�\�.9[���q=#��W@|3�;9s�*��۲��{9�;��������j��9�f:��]�V���v�&�k�;vZ��~n}�Q��۳�wa �J�LL_�����������V��n�_}�}�� ��)mZM�.�t��8���n��� ���s�5���F�	�T�(I�i�����`cu�b9������݁�O׀w���s武ݻn��c�vG�3��v�c��i�:��%�ə
�T�%U]>�w`lp��s%�����Oπ�=�+����v�6Ӷ��ո�i����ۋ��y:;c��Jy��	�������U�;�@;|��c�8��| ������ !⤦�եhvoZ��ʺϽ���Ӯ*9�x��0]�^�� �����o��ʟ���f:��"9ă�6gfaMQEL��S]� �ݮ��f;�yH������� ݴ����i�m;i]���}���� {v<�n��� ��T���Պ�t�p۱�Sv> wdx�vs�M-j*��Sn�.�v�ț9y^۩w���p槏;#m��;qv-m����v@� i�$�e+m�Sv> wdx�vs�ݏ �e*Sn�Mۻ�y�����s�ݏ �G���'�$3�Ut��N�$��7vNp��}�|�l�x����f�}�t.��OWhYb��,N#�����Ռ%06����ҥ�*D�]���Wz��i��$��n�s	I��t1��aHh�H�8X�`3b��P��:D�v*��� �>q\z��v�&�N�
�U]���{���w�	6<o���]�e7h�S���nǀuI#�vG���Q��s��R1�vեhv;�o �G�� ����=��lFÌp�O4�P���m���7 ⶟k��c����[&ס�nucQ��+Y&H��e�W$X����~�w[� �c����ryn�Հܤ��j��J��*Jf��fcwz�c{]�wv�ݑ�u*��m]X��J��ݏ �G��������'8��
U�*��
j����B��ݫ �ݮ��ۻ��s�8�k�{= d>TT��T��M�w�`cu�5r8����ok �G�;��ʻ�@4&|�ZcHI�ѷ�1��M�U�!أ;\\���;=�m���ͪ�U�b��1+o ݒs�ݏ �G�� ��w�`�Zt]*m�pَ����A�wv��v�cn�*F�ݵj�N�j��RH�ݑ��Np-�xݯT��t����;��M���}�ݑ��Np-�x��>�i%I�i�J�u�v�9��FN=���X�n�� S�*>�"y�"����8 mM��-(�0�R����Un}0��H9.2�r;V\K�qh���CJ[�;l4;��:���%�y���ns}��^��䓲�hI��b���߿�P�n��rnf�pջK�l��� �ݎ^�9��:��l������;e����)g/[O�:��$8�����훮K���'<� ��֎s6��笠��U���v�M�Y�b��H�U�+.۳��NBzV@�[���(���z�u��a����A.��:-�]����{v��1���ќv��g��/Qڤ�q�.�n�$%��息����mՀ}���DG �m݁� �M@��v�w�{�$� w�<ޛ9�<����PS�M�m[�vq�� }��{���DDr���{�m̀���H�b�QJU	MWC�!{5��-�� �od� w�<{e��.���:(�������s��X�u`y��7w~� �b��E|�q˶��5��.ۃy�J8��s������Y}�ĝtVy�;�<��V��uiݻ�8�����������X�z�3�0�k�RT��f{��Uߟ}�ivȌJ�  )�� 9Y���@yI/ �#��I(��V�4Ӷ��W@�3�^�=7����7�V�ݮ��A�K��J�I4�5v�ȎDFN=���ov��7]��w`{ 5��M�Hm�Ż#�}#�7۳���/ �t�*�O��wCo��rӸ���p��۝�\h�=+���j���׽�UCtVSݶ�ۺ�o ;���w`y{�#��A�׻V�ӲB���E)T%5]=���9���@�kݫ ���y�p{�u T�P)�w�������8E�*R�T*UR����e��������1���nڻ���&�� I6g ;�<I��mȰ�^�-KI[����-<��� W�U�ٳ8ۑ`ٳ>�ߞ����|��h�]���;A��]�vxݷU�h��fvŸ����u��e2cU��R�SIL�X���%���l� ��ڕ(�nՊ�t��p	�"�Ds� ���<n�ǎ�`R�b+M�BV� M�3�dxٳ�mȰ�PS�M�m[�|��gy�\��-{��3u��%���s����%2$t!YL@�FHA�
�� h�y���Q�PHg֛E�&ZbM��l� �UQ�uXz�� ���B9�H���Iӌu��uF۷!�I��s�Vp��;oO�Y�Ϙ%1r��%䩒q��컼�mȰvl� M���g8<���[i���N�۶�vl� M���g8ۑ`ez��V�t�Zy����@�x�͈�" �#��;������-Q�li�m+��	�g8�mt���K^�t�5=JTTԩ&f�)��Kk�j�Dk׽�_���_{��u�]��d�0��d��B���R}_}ݑ��������e�1Y8�kZ�.5cf݇�Й�miv�b��e�z��v���]���iɧm����'g��G���:�]�R�5�Wn�[�E�=�ej��Gf�X�l皛�����ZG -�������q�6{g�����-��m�)��sd�&D��BWpn^z^6�0Nj-r6k��N͸lr5��n9{�s//M����˻L.X+ �c��*��URC��k�~�w�n�qj�Gvl�v�g���%8N��J[��Bv֮/n \3�d���*�i	M.�f�}���@y����r,��ݩHvڷn�m�� Mn��D ��݀�[] ~x�`c�qP���v��ؕ��M���RK�	�8�#�=6_�.�wBT��m���m�@�>�cuЈ��n�y}�����Վ�&ۼ ��3��<o�� �^�d��-؛+m:����s+ut����mn�$����x�Ѭ����bt�ݙao���-<��� ��9�<���U|=6g ��B���ƚvһo ������W�EY�d� ���� �UK�*M�i�wmo��nz�x�g"" �n�����*aW%*���5=��BO5�lOߞ��9�շ��@nԤ�m[�|��g 7dx��� �^ o�>��$��Q1��	$T*G7���������;&䑔�,]8�J�Z`�RJ���1I5H���3BSU�3sv�&��<�����Ԍ׳�٘I%

&��M� ����{[����ݜ�9y|lwm�ݠl��� OM����|��H;��d�$`e*�'>�>�u�~ߦ {W��(���Ǒ�fp<�tx����f��9#���!�{��J6E�R��jJTJ�:�n�)��}�3�o����J������'Cu���{>�Kg�ë��7g�sj^Z7�m��GI���A�u�[��m���� 7۳8�8`�'8�j�@;��ܶ�w0}��pUUUI����96Np)���M�H��m[�|��g �G�d� �/ 7۳8�&��K-H�r[$�RI%G>߾�*�>��r��=��u_����Q���V'?s�}߿E�M\M�i��wv��= �f>��L�p��݁쟿����]��֘|��m�ӌ�l>63�N7[m��m�Z�+�E��!��ѥ9#SS��c큞t΁o�DG9�<���k�.�WV�.���O38�p�96Np)%������d������%l�9$��RK������7wfp��M�.4��mݶ��e�]��۞�ff>����-���̂�)���M�HV� 7wfp��[m݁�۞��>� �G  �" �`< <L"�|}]Ԕ����/W	pH#���xx�۹)�����4xs@:$=�N���}�ͫ"�%@�J`'��Aܡ��sX p�G���dP��lT�V ..��bgpp�禕^�9�`z��.�.�Cb.�4Z��p���A� �/��R/�pG�#���ޭsY���7��u�	��N��m�.�V�i�b�4�\�i�����&{e�R�5V��I�]�*�6�X���%�-�]�������|݋8�
�N��L\p��npF.p�l�vҢ�����ƪlt��j��:�Kn���cY�����"a�Zi�c#��ܮh�=�-��k�e����n9[�T����ed�m�$�Gu֝��rF��B�J�Ѷ�v3l�4�t��� �[����c��� �M�g�:���V�k��pdֻ[�u���0	�6jU{G���`K:��g������q�tetN�Ι�N�����v�6��غݵ���g.*��+�rygAl�9��W:��%�����Da`�/9ZtmUR\��0�g�NjN�P�N�[`A@:�N�;�3V崓hG66б�RhvY����9�]90�sl�'2�R�U=]-]m�@��S=��Ý�jB*7kK2=���6��Ԫzl�8�CxKh+j�C:��9W�u�Z���FX3p�nN�� ��u�����e$1���1v��:�N�r-Vn�Z^zIk���,[Qr�U����{��m�{�&�U��&ݰ#PccHUGZ��� �X����Ժ��U���kH��Cu�@yb�Dꪕ�����[)KjL���C��CA/`��-�+`}M�Wr .����S�,N��
r�oFJ�Y�6���6�un�.��kv��];V8��
��v᪨
2C�e9���U�|�{^�ݭ��-�N	��v�oNzOx���H皼j��ZW+ڒJ �%�K�2�Yej��P
�4��UUU��үEx@Y�v�{K���#Uy�w�nWB��`�}D�k�l�j��������d6�`�z�mH��n�u��q��.��K�� �󰲵P �^D �+`�V�����nK5`��É���+�x��^�U[0���.� 2��v흹�Y`&7lU:����AP�_�h�D����LN �l�M"�z��	���E�@�|���-浙�o&�rS�GZ�����l�Ŏ��]�۹��,����8ي{�:@ŕ1��8M\�����xՠG�²�k�P�c�4�A\�9����+��m�ܔk��,u���qݗv�gVZ��2֧��ؠH���F�v�r�`����|�?!�]�g���8��']i���Ys]�j����&���ݰ��RW#��$s�g=�)�����w������Nx���G5�uj��n��18�	ϟ]�HVqnR���IĕRM�k�ݹn\��]�|߲���w`y6����pĜ�&*U
f�3G@�ۻ��#��vz �큘�؈��G!�V�J��E$PL���1n��31���9ȈI��:ۻ�`ˆ:��EI!1P�������1�:�n�s��&��Sj��*�+��e���v8`������b���DZ�{���%ID�fKu<�.{�6û)�����4M1r�c�>�v���ɗN�Z�u�������ݻɷ= �f>�������Q6]ܗn�\$�p?��g�8�^�T��DGb",-�l�֝�7w��DG)#`TK�P[������� M��p��rl��RK�;�Q6�+I�m7mr�y����c�ɲs�yI/ 7۳8��uj]�cI�v��&���$� �n���� ��H��mtv�ꉳ�un���ܛG���/=��ᒽctk�������:��*���y6����1�'�-�w`)�$T�J�)���{1����i�>׻v�}��i�K�L�"fQP���9Ϊ�߷�ʺ�߾��^�Rd �1L1h���"�o>����	�L��hRQm�cm݌Jف���DD�׻vn֝67���� �H\iScn�ݻ.�8�p�7���x����Ӡ[���y!��%&�鞮ҩՎ���Ƅ
{�q�ؚ��PE�٤z�8XSyHM[y�]���ܶܖ`�vg ݎ&���0�M�JR�SJ�i\�W{`f:gw�kݻ7��`�vg ����T��;�Mـrl���������0��1)�"�R P���6"9Y���߾�Ϊ�߷���碸�a($����H �@ȇ����ު=󭟭K��4��� o�~� ��tx��r��=��L#�i$�͍Z۟f��q��E���#S�i�g[���oen�N)�d�1GlR)po����_�ɲs�z\� 7۳8�i%#n�n�d�)��[���9H͝����l��P��*lmݶ��e�� ��@3ُ�lG!&���kݻё�^|���v�����}�3�n��d� ��ݢ�@�bm[M�\��g 7dxUɲg �� o�fp������k��\�\Q�E,j���8t��u�rW m��]#Ͱ��:t�ٝyʝg�i%�m���ݶ�0�g��ݕq��46b�5խ�xC���ݓt��nŠ���C)�b����u�͡�Uշ���:۷'1U��qV��;�m�h;�=�9��.:$n�mZ�*`
����J��^�A���U���-�\��뇌 F�Ϭ��tkm[�&7'.��%�s�ԩ$�Mc���`���	�k��%ݡoj��l�6�� ���=�m�6^�䗧��f��o���������@3ُ��r���C���ىٞ��"
���3guv 3ُ��#�96Npy}��m$��*t���}�g 7dxf���r,�iq\�C��ؖ$�g 7dxf���-���AȄ<{��3%$���T��n�v���;6NpK�`�d� n��		[e_¤�Li;��ST�	v���<��ݹ���9ۛ��詭�&r:t�Rb�p;m7n˷��r, �l���ٲs�z��)��C�N�I[X���:П��Oʢ�u���o�u��ߺ�)%��(�R��ڶ���m�� n��M���Ix�ݙ�=%�Et�CE��o�96Np)%��vg 7dxk�K���MS�*M�XX��=��`��[����#������d
���(���E�؇eq�<ŝYԷh��4Ai�8�p'��'pF&��g�l��tx��`y�k�Z�Y.RC��ؖ$�3��<�d� �� o�fpz�Kn��6�uIL�tx��r�鼈���AȎA���ȹ!@��CE�0R(R�` ���m<���~�@w������ҧI�մݻ.�8G#�t=��`ct΁~m݁���L�&]�;i+�`��3�l�=$� �$��t��j�:Ln�u��u�z�ۅ����&5l�֏fS�wm���`C��T�<��i6����g ݎ��v�nv-����װ��j�TST�ـs�Np-���ݙ�=�� �BJ����J�)�]����@=���#��{3�_�w`˙2�;�ݪi�Nۼ ��fplp�9���uX2���10s�$g'0J����K&o�LϿ�|��%��N�3�{c�͒s�yl���ٜ��w���߃�ț��Y���=[j^
:�v�m�t7�@�&�[��������~���j �-�6��t�V������[%��vg ��ސ�ҧN�i�ݻ.�8�7= ��}�=���-���#!���|�ҡݧm"���L�plp��9Ȃ�v�[]�CpJUJiUM!L�K���v�q���m��`n�EH�L* ��M�v�q�������:�Ts��&5~~5Og]������|݃�'f����^4m���6�uy	{/-���K��Q��=��q�ج��ݴr����U���Բ���-�8�	�g`���|��pc�F-8{7<@t(+��m�t齏zGG�lA��Y3ۻMV��>��:ӹ.k,���+	8��ڢ�hv�K2��n�E��f�g���p-��E��ΆXwg'K����wwwu��ĒJ��k��M���Ʈj�[��.�۫ݹܥq�Wp���Yѥ�\��<j�ݏj�*�5]�>��ƺ�c�_�����v��l�Gr#Q��o ��س���G���on��N5�s������M]+-4�W��;�� �wg8��,�ٕ�{֒In�L���Cl��Ds��7�X���=�t̬:���J�;m�cv�|���`}���K:�V��w`\l8��%}7\Z��������65�ǅ�܉�H[�� ����ќ<��(un��ғQ�m��遝��s���}~Հwh�տ���ݻ�l���w��ƒ��T�I$��_"""#�E��o.�y-���c�wyN�U*g�je�������f�|��,�=�����:�c���_�l��[|�[���fV�צ���~��͙�U2Tʂ��it����#��9y��@�����ƺ�F5���+l'Igt�n`j�K��Ǳmm��<t�^v#ϨŰNܮq�
��xsrnG�p��s����{�l��=�I#u��m[m� �}��I�e��̬��L����f��J�[m�c�p���5��0�~ŇbJUv�BB�D1�8k�(�U	A�0DTMD�2ԑEd�FS�=���['���Ef�(�i{��ټ�Fh�d��\z9�wﺊےRLE��-�d���C(E�*5avy�aE�P@^�G[s��EY�X�g��eRDNT��Ȩ�
'�Å�w���a�
�&���aƓ��ǜ�9��]=����$����Ai6�F���0�DZ��M�v���zȏ5�BԚ4/��w���ލ��͞+�cz�T�����(,�|�/�)
����,p'"�	Z4��AVt��L0d��4�=l�8'g�X`�)	�5�5�#��kK&Å��8#bh6�OQSG���^�G�Nz �@h �p� �@[�QЁ�����Ǧ��9�7ƂA�t;��]T�6���@��g@���v����=(�k��M��vի|��0��\����~�}�b�8�{̒�{�v5��{f��7\s�� �=v��Hnힶ�ŧ���|�n�v&���e��f��g8,�=�c�lE���g@�݅�`��<e'J�� ջ/ �e`�z`��s�I&������������乀{�:�V��m�����j�2�Ҳݤ���dp�;�l� ��ߵ��_0c�1(��(
%������ji�����(E*V�i&�U*�����7cm���X��m� �}���>��V������ ߷I'�!ӊ�.5r]�s;��� �y��v�ݝ�9�i�m�[s<k���Y�T��m���Wv��5n��;�2�n�0��9�7ƂA�t;��6�}��9�@^z��}�w`b�9����G�5Ƣ%U*�U4�M\X�Z`�s��-W���L�wԄ���h(TE)�����c߬���y��CW���sv���S�UDU%5W`b�s�>�}��y��@��c�y�;��pV����p�\W"��H\=e��6��6k�E�^C�ζ��yu�jr��N8I6۷�Θu��r��J�������,e���l�v��d���b���.�!-�����;��m�]��Ѹ�c��uUϷ��"��8��v
5� '��\z3�.v���s���@��ޓq��|l�ٹ�&��Yѻz]��OR�$�v�d��&�����>|~��:r[)[ث��k;g�Fq����}8�v���8%��ˈvx�g�7<]����~v:�V｟�`b�s�����e��eӫ���dp�;�l� ջ/ ���=�I#V����0V�ｎ�Y�z~r#���w��>n��3vT��m���Wv��5n��;�2�n�0��9�7Ƃt�j��;i����X7^�{���e�ߚ�E���ⶤ�[V�.\�8�C;$��U�y�;u۴R��Ÿ�Z}wݻOk�Sjej�+�vG���p[���L�wɎ�5����r�����%U���| � ][ηֹW^}��y��@�nn��!HSĪ��Jj�����y��@��æ��c۰�͙�[�I����w�w�e`�z`��p{�L ��GğYMH�:�b��� �}��V��ٕ�s�Omc\�l�n�֮{>������#�	a�[����w|I�۵�;�����@w�?s�j���;�X7�Lf��J���m���v��5{e��̬����g8��N�MS�ݧm!��Uߞ�Õu��������Ǯs"9_�׷`j�s�>� y�T��Wv�\�\0w�9�5{e��̬}�B{j���-4ճ �}��y�9ǳ`{7{�Շ@�<�jk�*(� ��ם�8T��w�M�$oY5s�P8��j�q�\n9!�0�Y�F���ߣ��}�}&V��� �}�� �_Ep�i'V$:M[���+ ���w�����/ $����t��u+��ٮ{������L�����oi+T��Sl�;�l� �헀w�e`q|O�0�J��0�{E_�O:Sz`H\iS��V�ݵj�8�l���+ ���w���%��/��}3�au��ܣq�>��qf��\yB+h�oL���8�<�u�R`�?6������o��{�������7h�bn��-[�p�p�;�l� �헀w�eg䉻H��R��LL��V�۳�8�IxvL���6JQX4+�ݻ���p^���Xw�L���p�}.�m$�X��5n������w�߹�5�~�\B������{�a����e��l��f�l����PY9��'Om,6��]!u�k��䭎u\�Ѽ�vKr�㱟S���ݽr��� 	B#����q�9@v��ƻm�"�q���@q�gV���ÖS4G�]��x�#r\��.�)�d��@�����g��խ��
hڞ�;c=�pk�ڠ���Zaʴ��}��9��lԜ��ms�3�p�JU���pkz0�z���C�Q6t��a��lc65k�;f����F'���DE;e:ٲ:�wd� nd�a&Y$"�)ɋ�w����{g8�l��&V�ZIQ���bv�L� ｳ�W�^ݓ+ ���l�.4��M�m7mo���@��t��r8��)�ُn��BuwN�v������2�o��}�9�5{e��(ݢYI�lm�վW ���ݜ����l�X�T���r����h�v��V&�;q�X:�'mAm��rm���F�y��l!����
�T�M�݁���}��7��Z�S:��[3!O*f�*�f��sϾ�>Q6!�8��H�s���צ�{g8ؾRԶ�'H�N����&V��� ｳ�W�� ��!w�һC��]�pMp�;�l� ��/ �ɕ�s֒Tm�%j��Sـw�����^ݓ+ ���{w��ϰ�Z���A��X�ʸ!Ƿv鵜�ˍp��v�$I�I6�\Ž��S,���5zK�;�e`�=0��9�7�НB�ӡ]��n��2�����`�(ݢU��lm��.��0{��8m:�KK�IZT�O���`=2�����S�&Zi�f�{g8��Xd�Xw�LzJQU�J��mSm�o�}r,�L����{g8ݤUj�B"hk��(���n���C�ݳ�9K�5<Fۋ�$�ꋬ;�-���Ym$���:n��2�����%��QR�X�ҫ�t�3=��)��G!#3݀�wW@���9��h٩��u`���������M�r���t<�t�]%�������T��ls��!DDq�n�@���r���~ܬ?!�*|+Ͼ��絛|��uLt+�ۤ���&V��� ����W��UM%�R�+iڢk���p��v�uOl�s�L7c�]�R��9��ڻpj�N��M;cm�����`��s�j����UP�e`�R)�vҥ*�)��{��w�ȈHk7g�{v��g���$k݅�&�)䪢*�j���k7g�}���>�V�{��q9R�i]]*N���
��0}���%�﨩w,WiU�4w�XyL�c���c�x�U~�åz����������U_������,�-�.sq�@Q�����AT$T�n�w⨢���=��������������G�����YS������_�_����UJ�UUUc�����������uH**��������������TQU��g��n��s���_�}��5����	��	(� B�K*$�(�(J��*$ ��B�(��@�)�B��K*$ʉ2�D�� �*%*$�**�!�� D!HA�ЉB4
RPH�� L$2(!�B��� RB�2ą A!B4�R�!����� H�� � @$� H�� �@2#H�� B���!!H$! @�PR
�H!	B�� �J/�1 F@�@�$� �	d	@�!�%�"@�@�
"�B$�$F �BD$P��$� �&@�B% 	�!� �&�P��!DaA$% d	UaE� @�!R�@�A��� HFU!�%FR@��`%dBA�BaPBA� !	TRA� !	Aa@$	D�`HF � �fQ)���(F%Q� ��`	A�e�eDHFd�%P�dQ	F @�`@`Yd!�eBQ�ID!V�!Q�$F�dA�@F�aU@$AA� �`Q��HFFTHF ` 	A BQ�`	!B%F��B !@dTd(BE�	P�d �`FPP�		FI`B �dH@��i	H@�Q�@� ��@�BP%!!P%	@�	P V!P� F �TP TeEX�R  �	 F�Q
%R$ �	G?����TQUc�������xti����AQU�����c��#��9����W��������1EU�U_�̏��b�����њQUz#_���kg����5�����|;:QU�����TU_���FG������?�����
����}xj������ᗽ���g���;�8����ݙ��9�{�ߟ�TU_�o�.k���WW����w���?���PVI��\���6V` �����]5��  �/� H�� @ %B� >��J@ � r����(H)BT�*"��R�@� *�R���     QUE�(@UT \    F  �"�@b �>.g]S�^�<G�o{�I�����5q�������A�@O\��f� /[���wy � �:j��}<�ګ����OG{�n7{��g�槛q� $�    ) P(v� >}T���N��N%���L>��:P)��K @40 @ ΀&��b   	� @   t�(1  	  ��   � h��    d    �(�P��F&�;�>My�_{��u����=��U�{ܫ��X�κ��{�co� )��\O9��9��ݽ��O}��몸� =��k��j\�z.s���y�J� �#']���5粼����5��>> 
   � X� �uG퓋O<����Яp �{�V/�J��6q:J��B� >�>�\�箼ü <���ٷ�wJ���4��4�n����n{��7v�3�z��ӏ��OS����y=99t��z||*�@ 
( 
ah�y���Ͻ��Yt�9�帍���z�b��r{z��m���>�}����p��((�<m�x�ޚ� =z1;����\�w����� =8zX������bz��   ��B��R�P  �#$�M� Њ~=T�E1	�!���R��EH�� Њ���j��@ 4 DHI�JQ `�Li�^�~?r�����̠ݕ:����~M��M�л��(�*�@ES�J ���
 ���(�*� UN���#��D�(1"D�B) H����HC�6�ͱ���E`��$$�@���|��:�a\�$ ��H5������^h���������Q��:u`�"�b�V!C[���4Ú��[���l�>�Rc+ �+(J�[?aIg�_�.q����kB�� �)?f�C;�dj�)�T������Ee!MI.�R"M�B�X@!A�
i��U���uI�",�Թ�S�GLv�Z"{�ۑ���/���&5�n_ܦ���L)B5�Z�9����7��i	L!L>i.jl�8l�CF�6Y6��	��0ٶP�F��޵�^���Na�ɚBP�����{9�O�|A�<H�� XD���E���7#;9Ϧ�>a�]ӟ'H�'-d�1H�bivg&�VYbE��9�ֱ�
kAS�� �����1�
�����E���D��w�\��6
����6(��{���f]��~�$'E ���ѹ��"B\t���!#WI���,Ȳ\i��N�-���f01�e�,�i�D��p����o.2��
v��h��>�f014&�D�jc���J�n#�}fWA,�i`0��;5��E0�T����\�p���3Y�Æ�a��Ц�.�a�'�:v.�$a��c�g�f�|K�	s\ύ��ą#��G��kf�?�:�D.Mm�]�E��yT��]�����+mK����D.�9ɮs�jg�9��]_:��mr��W%D��ū�b4�7��)��*Sɮ�c'��Z�JT��'��a�\�oD�"�S�#+�B%�� �!T���;�
˩�D��1�4�H,i�,i��fd�Jԅ4	�	J�\ �s҈���_{=��t��?`ۍd���s�s�:�%'Q�ԬHP��L����꒣�gF�����*9(ުq͞��+(��n�"x��Ք��ur%�	�ڼ�|C�9��5�F�Ir2��B@pڐH�5�	kV��%g�X�$%`e����-�1��w��.c��� ���b�Ń%A�F �� @���
�M��Sl�����0!D�1Ѧ2D�SF�uz~�	�q!q�\~~��iw��I5ٚ�!5����"4B�(QB�ᨉ�;l���!mTU�+2�T�ı4ݮ�s�ڮ咔?���`c�J@�iCeqŔ�J�_�I�N����)$@�~�7���d
��"�.SU�_��;����>�	n�S�%���
��@1>�<�H�]�]#�#q!�@��D��v
bh�$�� D�2D, ��F�H��@)��Ԅ.!�,	
�z��c�x����� ��Bg3:��/��1`��>�a��5����B����l�Mk��ޖ+�3��6�ن���MD�Gi
��F�>8@�C��y�)�������^N5��\�1�)�1�E=w��VV�uR�H����A�fW��2\5(˳�~EYnAP� �IZ��%�A8�J�o�`E!��E�~9>3&�MKJm4�E(�J�;H��	��)�3dJJ����
�B�Ć�n�}��*D�vq>~F%4l��(���pO�a
f��8F$(r��k0��S��/U��㻚aHR��T���±�&�e`O���2�"`�B+i�J}P�9�!�T��i	64�nP�W	�1s�x]o9?�JB�6˚	u�$+�I��ވ��SE�����yN2�.ЫM�9�TZD)��S��z�+�I�8\e���� G�c "�JFB.:�w7��I��W�)�O� F&���>H8�����!Hi�տq��`�!u)�u��E�R"@�1?a\�4h`i�`XBR~iG ѳF��>��!.D�7�m]��n��D1D��I��%�%�\�$C���Q�]9�l.��5��XG4~�cP#P�SN�i����h?,����� ��x�`���k����>�b��8¤��B @�8�������r4!y+��3P�:a&�3�`HA�t���BRG!S	d"y
f�7[�:0���(B�||l۠�}:��#�"����m].�;��-Tw�˯�>�؛��5�2�kl.6� �z�H淏���3\ְ��"U ӓ'�k��$�sZ�7��t���K���$����S`ĬJ�������.�;Yx��$i�0��1�r�laXԁ�r��.j(A����	Lˍ�3�n&����Y�asIL�ώ�Ąs�k&R4�%��5���$���	G;�M���!$N�-�%`I5`A�!��Q�V�W��~-���;P�֮�n�|I�R`�1�q'�ϴff&�wz�p���te֌B��ee�K�(�Je��K��K��j!q�)*i�TH
jh�j���&�Ya"B\IV�5�]�6�Sq��]IL��-6�$HCX6�(�~~�a�1�e�)(E�\˒�C��@c�!C.���À@�2|�p8�~zXB7���@h�X�1q"&�ȵԐ�����v<�F'�T*��KD-�g9�Epi$c��g
K��_�i��sI�f��E
bcX���,�P���WJݮ>�(c&�g9�v�F�!qÌ��i����>b�!O���ϸϠl18�o5�������qM�t"W"��@@�k�^]Ή��$%	������,�J�E��NWF�~�}���]c¡�Y
ƱY���XBH1,+2��R4%�J�!F�HV�ꨀb�+��C�C�M�!Z語Y��x�G�,�� �95�K�Hٚ�~�F���8h>?	�jb�i��M�i�H��?��	
PLT�U�Mn�d7��O���H�3D�L4��<�jSH�� �:�!,#P`����D���FBH7T�Il-�`�$2$GG6N�\�2�Vv�:%�L%cB���>.a�ĶP��V$�#!Y͔���Ѕ����f�5�D�.�?0��r���[n�A	�<�x����6�Ǵ�UR���0UEJP[ ��S�'�?�"�8�o��>�рȡ�ď䈍t?3�JƓ_G0���)(���K��1�l
� a*K�ZX'�!>	_�{��h�i��8Y��j~����h1`A���?euHo�a��s��\����{�et�!W"@�A�L�ω�ˈ�T�B1r헭s�}H���Qգ�o�v�5����%r���k�j����(~�U�4�|F�FRc�		u5�d �"�ɍ�|��b�@�����%$G��W��Np��o�k|�D���51�A�q)��iF���5	J�H��ա(K0��k
G�P ��2�X��(d
���UcIu��V\��B*����}ϯ;�?��Múe�!CDa
c��V�ۚ��F�]:��!F%e4w��������M�2�KHRY��l#��T�A,JhY���V���H��b���B�UHP���bP��u
a.�M�M*y܅�5SYds����*�arg�*�o��/,џs���"��i]�X� ��Ė��C$�� Q�IR6%,BWwt���؅�~�ٲ}��) 0(�(i�]�?))u#el#��l�
as��tL%�[�Z×$�uλ�;��%O�YZF�H0,(B��%J�F��
��*YjJ��WI�J���G��������@C�l�X�A	 �� ��oY�Jܷ_��U>~�J�h%�LVWK��ka]xBM;�- T�����㤒\5$�m+.P֝��3@h6WQ�WN��2"�����̫�����n}�>���^���bD���B bR	��P�|�~ �L��%RCe��;J�]hQ-���y��	l� 	  �   H   -�  m��      �  tm�$�l 8      $ [F� �   8      ���       [@@       ��� �   J�[:7"�@ ��uÖ@�ג�)$"���.��!;W@�ĉ-�[u�X�p��ko��m�ٖ�PEm�*�X�T -�!�lH ��5UUJ��T,�>@�m� ���j��6�B\F�s�M�
M)�OUr��j�f��Z����J멕�C]�ڥZ���Io@\��mV��  l��t�s���m�� +J���^e�h�ng�e[j��5�-� ��M���m��]T�V��n5(8쪹f���9uIS��R�Ͷ-��ݰ����e��fx�'��R��Q���q�q>��m���Ӛձ-�85�`�4�ȳi�� ���=�q��ͣv�69�e{On[.��X*d�u�Q�Ȳ��:�[��B��Yy�h��,l<sQ���J%�{L;e;):��>UU~ꐥz�����]��q��i읝ۃ�j h�KUf�7T�eYy����� �!�"�NkwC I!��t� j�i
��dxа�N:�L�[Xjѱ=�8��:P.t�6�J���g[���G-�l��� l	'Z�#[�:X��#e���en�&��+�*�h3��é�k\�y��DtB��v�2��2�5g��f�[���@^�̫��UN��[L�]�l��r�   �t���n���  �p-rNض����M�ɒH H[C�ж� *��!5QW#������\ʼ��������5nʫ�* u�7U�-���k�MO��8q֒�h5�`��6����6Y����T�FY9�r�7e�H $ ��v��h8[mu��n�H �vppm� ���l 6�k�����R����#�*���ee�V���k�� ��-�  ���e��m& H���}����   'BY@�6غbM�R�[UUI����Zr�B@ �`�����YR --��/Q�lPva��`�ѳK�Zl�M�� %��K(lj@  -�h �]n-�l  	�pÃGP   �
�i^z� <���[U@Yv-��Iq�K=K&5��ض�I���$��@A����ΠA�ލ+ko`���/T����$m�  �
]��Z��jP6B���T�-��`�*�[qz�M���m�ְ  .Ki�oON��Ie���*FF��:� 9��qmx��a�e�����H2٥�ԆҮr�0�ņM�T�%�ݷ(ְVt�N�*5��MM�Z�v�i�`-����[e�<��"NLa�v�x�e�*]�ؔ0��0و:۠�
���"��ְnհH�ڬ�,�5Z��K"[;Bp���Ikq��&N�F��i�[*��U�W#� ��� 6���km�  �֎K(�ں�in�� �KV�m�C��[@ M͚�a8h낶�T
�u�J�V����������i8��&�B@�   6�Zm��j �ڭ�n�$ݶh�il�P�@�D�v�����Wnlml�pz�� ��`��lkZ��ͤ� �uHS�ʴm�����皬���IlbL�U*�HMUm�Z��4v�� � [\��6�m�m�ų]J�
�m۴���R�͵� �`�I}=�o��|�l���BtlʁCup�
�l�m $u��۶Ê�⪶Wvg��
۲�]��=�J�UR�0vx��ol�)k�i�`�]�Y猝��C����.�pq��\�*h��&�V�QOҠ`�k@7�*`�p�lkgJ�\�!�Y:ɀF�fY�� � 5�9�@�i' �齓P�`�ִƐm�	m�J��I%� h   �|}��@uO+uUcl@s�   8m�@��V��AyV-��	 H�m����� vͳl�[��[�N7�i$6�D1  �m&���H$p � �u��am�I�� #n�`�K;T�%�8����� ��8-�����   �u�i����ma��� �l��  � �6��	�Cm��)�٪��UJ�W�=�z�*m�����*�V�UU� ��[Uqi%��v�mR�k��S[T�+��@��	ڶt�*� ��-��Am �l-ż�l�8l�it�m�Hm� ��݆Vꀮ�UU����T �m�� 9m�Z p �d	�$��(WHL���U*�eقYd�Y0��H6�` m�[x$B���hkWM�[A��t�@H-��5ꏤ�pumD�(H�Vî ���� 	 l�ݶ[PN�`�1�iy.�  M��eN��Uݺ�Y-����j�  �M�m�����LUUP z�c�G#����Hr�,�Dغw9�΄3<��˽ln�Ƽ���b�B& �˳�m�u��O&3Jg1GJ����(6�b�h��r��mT9Uj^3��[T;����h�-��8Mkl��l@	      m<��b`�^[��m�k�* $6��XvK(  �mu�m�(��m4�`� ׭�fYD�-�nI+[ۛ[N魫Y�í��8 %�ր     -��L �� ��r�m�  l�l�`�m&� ln�'M�O����r,k	���� �` I����`���k �e�mz�� �ŶAl�m l�M]zt    m� �  6ۀ�d6 [M  6��/ZZ��`6�	$  r�����Ll'���x  m���m  8    e��� m��lߛ۽��m$K[l6ѫv�86� �U� p�gkkm����*ΠH K( �nn�6[�M��  �� �m�-�  m�۶��[n6݀  �   �6�I   $ $      �^�  YMkH 8Y`H  �2&�n��s�����    /Z [D���  l۶���`���hh     �x :sl  �ל p|�vp  l@m�� ���EV�7iW �smڝD�-��Z�kj۠A��
�T�bN��Z�k�In� �� ���v���O�|�2F�\sd��'j7=Mxtl[I����� ��D��Nm�4�m\��Nl�h�g�]�ȹ��D��j�$$6ۍ�U�%���U@@MSP�Ͱ  m�kukn� ��hm��     �^YYV��7I�U@W<ڶ H:��  �8� ۶��-��p �` ��i�m�+5J�O<�Uu�+��[N�    �6�  
�U�A�U�b�A*��8 �i%�K5i�� ��n{�����Z�PRʵ�jX�W*�@�ޠkm�>H��  6���ӧ q�,�]PU+r�U�E�ZVc�6��m�9�m��  {M�]8ӤM�9�[M�� �hm�[�-�Ӏ��m�l����lm� $��@�{m[6���6�"L� -�-�Lp���@$��e��	 �)m��^v?��o�d	��ye�l̼�g /KT��nͲ4ɖ�$��d��m����܎�:dn�� u۷ee]v-�we�`�-`�m�5�--n*L�V����P;'i�Uq�e�vv^�FԤ��:l��YEv^����H.�9�׭���-��v�� p[@ [@�I�q�=�ki7�����޻vض� h�m� �&�sm�lI��pm���  � �m��[�s��M�]�6̀p$v��Z� �jݱ���m��V�bθ�	�"�p ��2� ���tV�e�J��b�`kmjC�T� h�m���ݒ-��$�H\��WVÓ�ۤ�c�����E�ݙ)>Ҥ]0l��ٻS�����N�ɗM�� [N��� ��[SӜ��6���N �� �m���UUyV��ve�zUuL[��f���; �k}�8݃�@MM,W2�T��giUmV@�`D��Tə�����FKH;W*�O5^Ӣz�ԡ�V�r�vG������*W�С�lfU����|�kğ"�T�T��i��[l-���� �K�m� �)�K( ���붥m���m�p ����~/��I�8 m� m���lZl�U�� E)�� Àm��q��m��E    �زҸm� m�6��e�	V��z�*�i	T�ہ��T
�����T�@kUn[� 6�ѵ��Ԛ�!)�&��*����Ā�����������_õǈ@S�"�|��[� ��!���0D  "�7�(D
�Aq   	@�������"Qئ4����S�!ޏ�UA��6�(P@�� ��4�t�����	�>��X����UM ��Q^�+�<E t? PR��O���q��E������� c���E�� ������ I�
��B(����>�(T �x��P���#1CO��D�A��B�Th�	Q���#�PS�X#��6��D��*���:�;@�pS�������!�PqD>_�A6��E8鈟�GI�>Q�^�ׇ��?�S���C���]��!�h4O�P�DL ç�z�T�5��w�H ����� �"���єN?�|�HL������0�D���L�_�Ƒ�"0Ҕ����A~��E"��0q�^��ʪt��ߪ��A]� �N���.��/u��� �a�������QS��EWj?��	��	D�Ab	b,QJ�B�E,�`�@�V ��E�Q@��_hֵm6�l�m�� ��m7am-Mxlt� �[v�K3UGΫ%�3�� k(N�+R��!��bG�t^<��}����"yN���j�ўS�)
�2�F'άvv]le�u�.qR�����}�[m�wA�ɚ���z�!EմIu�z��]tre�8k����8Է0QjR�eS-c��̭y��Ύ=#gk�h
�Un����c����Gc��ji2��uh
����a��e`�:&��TP)�jZ�eZ��Yx�a�ݓm�6�C4��OK�Z���ͯb��Cүt
�@��Pj��c����EX{��S���'\��cLv���9z^�<]Z�Ҁ3�ںx�M����EIВHS5N�8�kH: �v����72�%�+�(T�R��s�S�ۻI�"}��0W;r��`�N����n���G==�m����#��E�᱙��*�A��vmY]�n3�;�.)�^Z��4�r�ˮj$�HY������VC
ˍ��lWln�{��{c��2�/N�u��ƍm��a�m=tp��
��Zr���.��n3�eyv�"��];۩�1������B@��V�C ^�A��M�bԳ[���6�]3>L����⒩y���nX-�]���yBv(6���]�zngꝇ2��\�C�-s��H�ZAm�-�A��u�I��M� 5��6� ����-�!�;�u�˭�>Lci;e��u�etk��Rŕn� #]�2����I�.L5J��X�3�ۚ��孪G��;�r��8z��ͭ֔���0u��
�)�0��T�{Wj�ʚ��*\��2�7Ah����
�;u4P;%�h��k�	Rt��&gi��������C��I��9�V��ú���H]��'e\��WۖӀ-�t�qٮv)����wa�jj��wf��Qͻ�v����m�^])&�Ա �qWzʿ(�u"t�i�L�q�Db!"	���i@x `q�N�>W�
�}�~pa�^v�O)�e����t�k���S�]p�x�$V^֭�c���bS�Ta.��x�M��-�=O-���	�ҽ��:!u\�#��\���s�c�hL�!��s�������ۜB����fТD%Wg u�*5�v����6j���ǥf����_l�Rn�v���E�ݹH�V[��k�w;B�����F�+�^������^�y�F��ݑ2<g"�7��¸ۗ�8y�x�3��c��P�飣36Ձ��(̬E���ٰ9�80���$��I"iXܭ/�OD�s'��(�"뗠6�ց��;��]�,.�,W�����F���w�JI6�	א�;/U�(,@�A����@�ޯ@����Қl�h�q�X�����m��=�)�[e�@��w�IQ��E�e�Ve	]�P�8��q>�ZA2s�;97FK��{J��Bb^��bLk#�����\4^��m��;�w°!#	17wkQt�+�Դy�T M��vLg�z׾��=�)�Z�6ٗ���+ř�h_7zm�i).ǐ�$�(�<���YX���8�@����;C@�d�@����?:���bN��HB	��=�)�[e�@��@����\X
~f\x�,o"A1�z�.ȴ�A�۝�]��+\�u�y��Q�:Kt��drC@�ˆ���^�m����4��\�$ P�����C���^�$�Zϸ������
8E���m`ۏ@����Қy���ʃT�Z?#,�@�HhoZ|�l�,�ݛ;�+b���b���hޔ�/;qh������<��l*h �	17����^�z���ҚT(aP�k��$���g�6���ݴJF�z0i� Ŕ�ƹ�w��W*�vmU��o��נ^�s@����yۋ@�Sh�I��BGz�w7��ύ������^��ǔƘ�cRHA���>}�h��-%q&�%�ɵ�~���27���G$4��Z/m{�w�{�rc�����i��59UY�4#�ŗ�ZV�^R�2;�6�������;�,4��w���O��p��կA6��#��z�;^t�F�M	֢E���-ml��Uۊ`ˌ��E���96��q��Js��U�|���)�$�c"��s4oJh���^����i�<��x�0�p�/;qh����__���;�>4C��2���Q�$��'8��K��k@���|�Z��Sh�I��BGzu��������ߎ��yE���ٰ�\iڴ�R���([t�Ȩ��])X �@LD��"��P�D�	��b�1J411Pp 0��C��ݟK�a�.	q�W�6y)ݱt�C�Zn�S�m�F��b+����X)^�Mcm�t@��W��ΰ�8ѭ���3�n]Ѷ�#��n��y�=��!�e�.&��a[7v�g3V[�=үq���-�VҰR����n57j�Ȃ)΍��q�k�xq�e��k`ڮ���YKi8휷�C|o�N����d��B�qi6f�Ճ1����� ,16(c�]�ƭ�8P��c��_'U�YC�dq6{+d!"�5�16%Ӓ�I�~�|h����^��빠y�do0U�E�y�h�ۥ�W��엠v9��{zS@��{�HP#i9�@��@����=�)�w��Z+nB�Y�fd�ɐ���ܘB	КBc�����綼X��Q`dwu���u
D�8a1�3@����߭�ZW�ށ����%W'ej�
 <��i�5צ��y�.W��˼�g�D�q�;c����vKb��Ѯ�gj2������R����>}{R����#y�c�HcɍErI�@��^�~����d4�Z�P����V3+K;;�,)�<U16��H�@����/t����W���rf&�\h�a�
�%W9�Q����rR����=�w4=�3L��员�RHh�n��9R���6����;M�߁�qgup��78��Mv�6�r�ٴ��7����<N�Obm\� v�(3�W����s@�Қz�ŠUԸ��$6(�`ӏ@���߿~��96�ے���[� :V[�K1*SB)L�+svՁ���CV��ٖ���Z��f&�6fm��m"T���H��4�ۋ@���o]��w4(c����c�Q�&-���޻��w4�ۋ@�w��&� ��\2�K���p7����NS7k� 1ڭ�����g"�,*�Ԕ���?:�h���;�n-�k�/�&bm	�ffa�
����UI�%-'%�>����>r+4���*�)ZD�4��hu�@����/[��yN�Z��	���Nb�*�^���rN��vnN��8PV�����z�y�-�x����lQ��������$r~��>ܔ����|4�1�-�#썼�(�M�Rn��jCvn�O����\,�(9c������h��WZ�o]��K0�+`�Q4�UEER�3�����I�I	6�nd�z�6{}j��ݵ`sJ�,vO�����LZ]k�=�)�^�s@�]��T�I�	��	��޻��w49ۋ@��z{rf&�+�$��	��/[��y��Z]k�=��g�. �i25�ۗ9��MՕ�"m����k����r���t��>��������:�M�K�~]�k�����q� a�M���^65<>��m�����m�vӰA���LÝk`{��t�v�tn1�ѥ��g8�e8�W�X�`�M��D]���"mŇj����'�k�ݝ
�Sm瘵������#Z��6]��Rq�Va;hc�z��n:�f����]���o����z�S<���v��-�!絮��-�T\'m�XӋ��Fch$��{���ŠUֽ�빠^�s@��&�� �i�Z]k�=�)�y��Z]J��4�1�6��=�q�)/��K@��^�w�J�ٖ�F7D7!�^�M�v��*�סqu�s@�0x�aH��s'uE��KӞ�����s+K
���U�9##�Pi���A�I�(���ط>�W��۫��Q�b5�`�0rs6��V��I��J��z�K���y�I^�Q��������������E��aNY��Lݷ�g{�|s�� @���$"�a
6�J�ӥ�]]w^�jI.�[��J��z�K�����+�$��	��Ē�.�RIy��^x�Ut�ԒW��<�$�t�_��~Y1����$�Kqy�IUҏRI^���Ē�.�RI[ʴ��@��s�s�$�](�$��K|�<I+��5$��n/<J� �}���el։%a5��˚�SS�Y㋘ŧ��<��v6��>���-Bl�D#��$��}�y�I^�Q�$�Kqy�IUҏRI.��n��d���y������wf���������[o�u��%�_��<�$��L<�@��&�F���-��$^�����30ϖ/�3�T�!���IQH	��3�p٥��,x*|Z��� Ȱ"��a$�Dd$1�P�ʇ�O~����{���z�G�(wG(?r~~����APیHFF@�
��o�HKl#YR�-RH1�ܤ$��M�xM�h{[U{X��M�#�u��w�֩��jJH2���9�x��hF� Jit
p�y�168����N*|���B��pU�>O�>*� `D��l.�g�9TҪ�U�SZ�\���9m������m�J�V:�����L^x�E�I�$�[�_�$��=F��*���=����%�lF��7N8MI%z�3�K�]�v�{�]�y�m���˻m�3��?{��k��^�c���a͸�#����o�猾�
c$��7=�J�g����}�ԒW����$�ғRI^���Ē�ҽ�a�df6�F���-��eUݣ�!��J9?W��%���o陉I�_�D	�`�Nb�Ē;��5$��|�<I.�u�J���$�V(��1�$���5%[]o��%z]F����w��-�ѯ�%mTk�Fֵb|��Ү""#sL�LԊ��hW���IH�~G�_r=���$>�3RIw����]ݚ�T#M�x71M\������heے�gk�����JX#2�9v" D�"�R#RIw��/<I"��ԒW��<�$�K�ԒV�a�V,_�HE$�b�Ē/JMI%z�3�J���I%z[��>��\��x��!����RI}~���Ē�Q�$�Kqy�I�I�$��?"�*N)���%�.�RI^���Ē=��RI^���Ē��^�Ѱ��cC�#RI^���Ē��{��J9?T��IG�Q�$�UmUW�y������H+�ff�3��\v�½��5�i�%l�1�"�y�0��[��j�l�`��z����s=S��e���t<G���߫����=��TY��"c3u���!��{Q�ke�X����kd�Ό�v�\5�<���Г�u�lf���/r�(jŜŰ�;K�Q�/W�\��v�He����&M"�K�YZ9�n%)n�w��}ޏ���v��/�V�Gj�<� �]���������9��Nn۞v�d������lnn��ǜ�E�|MI%z�3�K�]F���-��%U�Iɍ�7��ۄԒW��<�$���jI+��^x�G�RjI%���w$M�I<M��Ē�Q�$�ct�~^�]�ِ�I%���$�̶
��@��&�F��󥸼�|�;��5$�[�x�]��5$����b�I$���$�l�Ԓ_��|��Ԓ�}�Ԓ^t��$�g" ��E#J9�b:!�E��%#7XLb�r<N�ccY�8�����s3^ō�OaO�''�$����Ē�q�5$/���z���;�I'��-I%��?#��_��r)�
C�K��Ū����r�W*֤�>���$��ɋRI}��7�����uG��������r��� ��|����;��\GͥHM'UY�~:��e%k�qjI/~ʾ<��cS$�Ē^�bԒ]n��K��ũ$�[�y�IWaRr0��Icmȵ$�[��Ē�wqjI%��x��ғRIy�����Y��p]�9��g����nPM���v���.%0;���R�r�!p�BΫY��Ē�.�RI.�,�Ē=��RIu�O<I/h�'��N2(5"5$��r�<I"��jI.�i�J���I%�*�G\1c	0�M�y�I�&�m�����-N H� 03�𪘙�g�'���5$���'�$������q�#�Ԓ]{i�%z]ũ$�[f~���/�6ZԒ_v���V�%�x��/0��$��{KRIz���O{�w�$���։%׶�x�_߭>ũ7��c��1�M�x絢��Q�`{knvJ����vyݤ�A�5��-���M�r���� ~���������$����\��I7�Q�$�u�I�D	���'�$���=������H����$���F��]m�����9ʫ�Q}�r ��Ibm��I+�ߏ<I.�=F�+��9ʻ��~��]S!z�I?�1\�6�#����ė߳�fc�~���{�zk��߯uٛ��
����-b!�
�?��Р߁�P-�����[o}3�\&�ԑ8ȠԈԒK���Ē��s�~�$��~<�$���jI/�S�<�g4��LݻO%��e����L�me=�!�;rq����f�k�,� H7&O}I.O�Ԓ]{i�%�.�RI.�ry�I{Z �'f
	�q�Ԓ]{i�ْٟb�=�ԒJzz����[j�r��/�Y�|�(�&,��$���F��]z�~��]�UȯRI8��$�����Z8�cC�#R_cn�~��%���z�K�u��$���?{�jI/9뺴~�
��������[j�$��ʪ�'��;Ԓ�=�ԒK�����|W� ��Z,�\0���Z��՝�ue�G�y�m��\a�Z)�v��Z�uZ�=DV |��F��f^6�i�3�u��uGiTk
�C�/K���Q�s��T��5�k���i{�I�g�}��;ΰ�H�Uَ*��-��.�@œuU*�«���S�>k�199��ݧBY�s�WX�
�wdxқ$ͮ;�UŞ�[J�7�4h�%@|���[��Z��r^���2��]]�4�y:����x6:�s���N�}����h������7���%���jI%�ْ���]W"�I$���_d���4܇�$�t�����m|�M)��}�Vl��X�ZXqh'��N2(5"���@��)��W�>4�~Z��"�H�c	A�	�y�hzS@���h}�_���}Q��	D�A�4�)�J�q����?|���h�����<�跭��qۉs�vX�ל<=Wv{�6�����Go��|i��`�k��o��~Z��h{e4�)�x���q@�R�f	����Ү�	�]JM֊#.]ij��~ɿ��M�ŭ���ֶq"t���n T������3@��!�u�����]�s�@'��4�����WVZ�"��xhN'�@�mŠm�����N�\��ř������a�}���޹�xπ�-�Jh��S�`�Ec�bq,MN�z��^�*N<�0�m�N���>v�-�>���a�Q����XZ�_��)�x��~_vL��!�s��n-�EX�W�YH3+(����ͫ�&�NRK��Q�_]�- �l͜����.����X+�%EUU����`s��KI,+��JRI��k�O�|U�w}�X��+TIWfe*/0М�_wZ �h��Br��a�|���RV�eYv�e�����')}�3�<�����Zi�7���ŝ��k����%����h���ٴ��7
'k1l�x�ڟ�w��Н�lq�$<m̞ {��u�M�]��������-�&�1��F!�&�ץ6r�>�ȴ����͜�A�j\�$Q� �����z��i���Wcs٠OL�~��+��eb��2�+�ЕĜ�� �\�����.ꪠ��& Pŀ@�B+! V�b���~�ZB��H.���;����=�V�dX�J4�3@>��4	T��~�܋@:�3@��g���];��6��5��iڷ\d���u�e@�fַ�8��g�}��y��E���Y���q�4�[k@:�3��U}`7=�]_�]z���WF^ﭵ�K�sa�޹�_q�)#�ڲ���YV]�Yx����u枯r�zg��疀����[�"�b.��Ћ��@q�4�_Z��8���>̊�39��1%�b�Z_q��wv�p}�`s'6,��i�&�� 銆�������O�������,	"�$B#$"H�"H,�AtQt�XP���H�(w/�t�_�c�9'8̼��y�XFA#��4��#LH�;� �ຄ `��F�||��J˳F�!]�`@��B$"�dRF��1bF`DCc�iP��ȯ_g�.$e�\h�Wb����Z��삆�"1����!� ���!1!�H��~ �O��˿��gn�Q?,X�4$��]���®$�4�Ni!,� �! HB�'v����vy��޸���<�C�[M� H&�8-�k5� ��� 8�*զ�K�	�����n��*���ڧ�^pg�Kb�S�l8�y{Y�|cp�ɽ�]�N
��J���D�F���ol<We�Sf������c�N9���҂��p��BT�`��!�l���Aƍ�r�Z-�F;i%���܋!�\F���Փ��3iᑫ�:OcMm�W)�z�֮ݎ���W=I���C!4�� Q@t�J�c�����uI5�d.z���`�l��bu\���l��\��,���p���� c.c�qN�<�� N'�n���92���I�i%�eg��˺��z]��l]�ɰ	n�kH���`IP�〔mY�]pl�E�[n��ix�%�z�=�˥��U
��5���e�:�|q��l�6�����e���jxSk���U�+ֆ��Vɺ���v��'�Gn�]U����#��Z-͍���;ح�N��uR�M����[[n4�ʎ0��[m)�F�����NG8re��\��x5��ƣ����qu�o6�+���"�*$g�}Y�m^9^�Վ�-'�"�۶ y��[�[�bn��^�CM7K�i�vYZ�ck�V�,�nӔ�0��/[�ٽ�h�2`��925:�6��$��M /P��c��73�N�f�� ުÆN:ݥeC�e�`��yv�4�.م�ڠ�Z�7;�h�jU�B{m�˱ok�;N���[k��1�s��!z�
��!R��6��ҳ���ič�4@����!.��Hɦ`l5@J���dۇ,��LE�.Ԙ�ـ�'g��1Y��	��UV٨�^W�p���8��4.�)u�r�X�TQ�s�۬��pk�N�vNv�,�X�@�5m	�9�Ul�x۷K�n�^�gmC�WNQ�n����)��/p�nQ6�gl��lU������+p=�������6m���
͹��۴��
�t��[t䱠����YP6��I��4a0�!�FyV��������|i�� x�!�#�$?N����~W����P�КR�ID�PI2d�K��U#��w���Cű^���2t�m�)5Dw/M�su���.�cYs	�u�h�ў�j�Թ�3�ӌ3��@�y��k��8s:�z]J�w9[���C�,�;u���G�`��t��(݂�Um!�P���9v�쉻8�oZ3��勗Lo����
��:!�nF�2U/7X����A�uK߿7�wܭqշ����{���i~�V��V<�J=�M۶������q�'g��p�d/&����cs6�!�}�|h[I�yϪ�:����Z�o�9����4��7�Uď���C@���4�XGT�a!m7	�yϪ�:������U%�y rC'*�_�6х���"�<�QH����Қֳ4?��-���R�Z��)Qw�����h��������4�W�����~p��v���r��혠�v$���5����4�v��cb}���`w�ڱf����o�i8�R9N=��0>��,K�����Kı?��JsVJ\����jkiȖ%�b}�w�i�QҤT�>��#I*��X�idMı=�o�iȖ%�b~�w��Kı/}�Mm9���2%���o��ִ㚚��e����Kı=���M�"X�%��{�M�"X!bX�������bX�'��}v�������USP4�&d����K���~�ND�,K����ӑ,K����ӑ,K�!�^�����5P5Y�	�t�&����fjm9ı,K�{�[ND�,KO����9ı,N����r%�bX�w���r%�bX�=;��r�W&:{Bdz��g��F�٣]��n����Q��݇9��F�v	~�wxS��Y��@���9ı,O����9ı,N����r%�bX�w���(@C��G)O{�o+��G)�r�����-`��˫�]�"X�%��w~�NA@�,K��~�ND�,K����ӑ,K����ӑ?��"X��i�Ҧ>D��f�k�P5P5���m9ı,K�{�[ND��~5Dȟ����9ı,N����r%�bX�g�ܞ��SFL˒涜�bY���"g�������bX�'�k��iȖ%�bw�ߦӑ,K!lO��i7�O�N��7P�aPJ��*�@����Չ�^�1S���6��bX�'�ﹴ�Kı/}�Mm9ı,O��y?n���Y�I�vp��t��1ώ��cE�x�W���}�O�٪���2}��o%�bw�ߦӑ,K��}�m9ı,K�{�[ND�,K��{6����w��������a��K�K��{��,K�����6��X�%�{�zkiȖ%�b_w��ӑ,K�﻿M�"�%�b}��˅�4j挚�jf���Kı/}�Mm9ı,K����r%�bX��w��Kı=�{�N@�@׳Ћ�E
eTTELL�V��bY�"g������Kı=���M�"X�%�����r%�`xE 1�#�sE���F$�UĨ���mSb��~�"���}��5��Kģ[��d�#�&*"U�j����@�D﻿M�"X�%�������O�X�%�}���5��Kı=���iȖ!�����v7�����F��.����a͌;�<�<�^�9�n7�C'7no���?r[2歓Y���Kı=���iȖ%�b^�ޚ�r%�bX���ٴ�Kı;���iȖ%�b}����nFD����fӑ,KĽ�|ki�6%�b{;�fӑ,K�﻿M�"X�%��｛ND�,K��޷j�K��Va��5��Kı=���iȖ%�bw�ߦӑ,K��w�ͧ"X�%�{���ӑ,K��u�ڙ��sF�m�fk6��bX�'}��m9ı,Og}��r%�bX���m9ı,O����9ı,O���k3*��)B��&���5P5[9��k�P5P/���{�V�F�j�k>�}v��bX�'}��m9ı,H &� pC�{?˙o�횒�H\��k��肧��m���F�Iy���(�{�\��6.7�N���g�X�6�wMu��'nj�������-W� R�qsK].��#Y��;Ѷwb��e絎^� �N�7f[8�:��hc҇���ن`ݵ�����;skX�v��v�zٞ�g�*:�8�=�e^��k�N7a5H:�f���73A�C�����nN+u�7���{ǯ�;}W��Z13�pA��"�����"ëg���ܝm�F����#�iѫ�2kY�sY��Kı/���kiȖ%�b}�w�iȖ%�bw�ߦ��7�Q,K��fӑ,K����?E
eUD*���V��j�g��}v���ș�����6��bX�'���ͧ"X�%�{���ӑ,J5^���e��j&J$*jm�@�D�;���iȖ%�bw?wٴ�Kı?g}�kiȖ%�b}��iȖ%�b~1�=�g��ܹ�um�M�"X�%����fӑ,K�������"X�%��{�ͧ"X���w~�ND�,K���z�atI�M\�m9ā���z����@��5/�}6�	bX�'�}���Kı;����r%�bX�=җfId%�]Mu.��ۜ���ɚ����c�}��Ev�	۝�l9#ܙ��@B�B*	�����F�j�k'�}6�D�,K���6��bX�'s�}�ND�,K�w�ֶ��bX�'{���k4�5m,Ժ�m9ı,N����r��U\wq,N�9��r%�bX�������Kı>�wٴ�O�O{�Os���-���Y���L���"X�%��￳iȖ%�b~����ӑ,K��=�fӑ,K�﻿M�"X�%��wĸI�F�5sR�iȖ%��dK�����"X�%����]�"X�%��w~�ND�,	�S#^���mpj�j�ߡ'�
e��T5��fӑ,K����ӑ,K�����iȖ%�bw?wٴ�KģY�����5P5[�=�*��7#v����&冷�cPk�'^(p[����3t�zcP�Ά>�7���x�?w���r%�bX����m9ı,Oߵ�k6��bX�'��}v��bX�'�Od��,��5n[sSiȖ%�b_�{��rȉ��,N�^��m9ı,N�^��ND�,K�{�M�"X�%���{�?�nB�����k\O�X�%�����ͧ"X�%������K��)!��O�ș�{�M�"X�%�~����Kı?~;�0欔������kWiȖ%�X��k��ND�,K�{�M�"X�%��~��iȖ%��*�
�D�}��]�"X�%������˚�s�5n�v��bX�'��~�ND�,K>���m9ı,O�ww�iȖ%�b~����9ı,O��綾��ujd0պ���\���%i4�n^��s�DC���!̳���a�Ӎ���p5����{��7��������r%�bX�w]=v��bX�'�����Kı>�w��Kı;���	8h�3FMk	sY��Kı>�z�9�,K��w�iȖ%�b}���iȖ%�b}����r	bX�'�z�f{Xf0֍SZ���iȖ%�b~����9ı,O���6��b%��~��iȖ%�b}�w��9�@�u{���Jj���(��j-�@������iȖ%�b}����r%�bX�w]=v��bX �睏�Q8���~�ND�,K�=��3�Ys.jܶ�ӑ,K��=�fӑ,K�����r%�bX�����9P5Y�~-�@�@��>>P�w���<��ۮ3͢�^�������{=���s�K�0��Q�����n�&�~�}ı,O�׏��Kı;�]��r%�bX�w����bX�'���6��bX�'�ǽnՒ�]Y�.�]�"X�%����Ӑı>�w��Kı>�wٴ�Kı>�z�9ı,Ow^=r桎a��]K�]�"X�%��{�M�"X�%��{�ͧ"X�"�ș�����9ı,Ow^��ND�,K�{ޗY�Jf]��nkSiȖ%�b}��iȖ%�b}�t��r%�bX�����9ı,O���m9ı,N�ޓ2I�F��sZ���m9ı,O����ND�,K���M�"X�%��{�M�"X�%��{�ͧ"X�%��T�����ݿx1����w)�ȽJ莇:k)���}%s�Kwӭ�� �KďKk�"�h��`,�rܗH;�pu99A�e�C�ZA�Mc+;������� c'��%�ڽk�q���|���XՎщ����zA�3��n�(ܮlɲ��^Q��ȺxtG9:���x\�6���ն��š�{[��^=m].{\���\і3�{O\s�Ϋ�����{������n��g���V[�:�{v����r�r7�;�����v݋knO����>�3㫵���ND�,K�����r%�bX�w���r%�bX�g����%�bX���趸5P5]�ءz��b��(��f�ӑ,K���ߦӐlK��?{ٴ�Kı>�z�9ı,O߻�M�"X�%���d��,��Z�-����Kı>���m9ı,O����ND�lK����iȖ%�b}���iȖ%�b{��OB\�-Յ�5��m9ı,O����ND�,K����iȖ%�b}���iȖ%��ȟ�����r%�bX����n�e,0��&\�v��bX�'��ߦӑ,K�����iȖ%�b_�{��r%�bX�w^�v��bX�'�����wFC��r�-�qWc���<�vys؀�lqXN�a�3�����mǗ�����N'�,KĽ�����Kı/߽�m9ı,O�w~˰yı,LͿ��j�k��/A4�f)B*�\ֵ��Kı>���m9GpD 1@�F�M%E'P���|�&����iȖ%�bw�w��Kı/����r(ؖ%����d*U
i�56��j�k���k�P5P5�������6�ș����ӑ,K�����ͧ"X�%������ja�5�jh�3Y��Kı?w���r%�bX������Kı>��ٴ�K��׳ٴ�Kı>����5sY��e�jm9ı,K����r%�bX��w�ͧ"X�%������r%�bX����m9ı,O��!|d'2L3V]jP̹�nw���l���x��ӮL�q�'E�6sIs�m��ݸ��g� �Q�����7���{����ٴ�Kı;�{=�ND�,K�{�M���>��,K�����r%�bX��ײ�B\�-Յ�5��m9ı,N�^�fӑ,K�����iȖ%�b^���ӑ,K��;�fӐ[ı;���d�[-�Vf�u�ͧ"X�%��{�M�"X�%�{�{[ND��{i��x#��lʚ�/��A���"Mif�HK�u�6��9�>X�5��P�
���̡�,E�s�H���>��
m@��&�c��q BF)"��,�t�詪h�"X@�K"j2ͅ ��
C1�+ �	[�w8�����U>�A���dA� ���H���T���t�6Yo���Y��jb"�����<z��"��(��z��*pO��z�����4���"::	�z��� z� ^"T�D�Oٿ�ͧ"X�%��u��m9ı,O{]=fkMs�5��M�"X�%��k޻ND�,K��}�ND�,K�u��m9ı,O���m9ı,O�~��3T�L�	���Z�ND�,K��}�ND�,K ��{=�ND�,K��~�ND����2'����v��bX�'�=��JK>�lr�3gS�l�{]�9�n�Qng�*�ns� �g>M�׎ݴ��/dIM��~��,� dN����ND�,K����ӑ,K���]�"X�%����]�"X�%��v���ja�5�jh�3Y��Kı;����r%�bX�����Kı>�wٴ�Kı?w^�fӑ,K�ｸf���e�K�����Kı;�o�iȖ%�b}��iȖ%�b~ͧ"X�%���ߦӑ,K�����=�ɖ�Ve�56��bX�'���6��bX�'}��ND�,K���M�"X���26�ﵿM�"X�%��wyBfR����չ�m9ı,N�^=v��bX�'w~�ND�,K�׽v��bX�%������bX�'�O���j]���훳*p���=�����iH��N��=���Ϟ��P�r0`��eK��w�{�K���ND�,K�׽v��bX�%��m9ı,N�^=v��bX�'����5�����Iu�ND�,K�׽v��bX�%��m9ı,N�^=v��bX�'}�p�r%�bX�����f�L��ueֵv��bX�%��m9ı,N�^=v��bX�'}�p�r%�bX�����Kı=ޞ3!8h�5�54Mf���Kı;�x��r%�bX���p�r%�bX�����Kı/�w��r%�bX��i���\1��MML�5v��bX�'{�6��bX��o���>�bX�'�{�ٴ�Kı;�x��r%�bX���x���8�aP�&"V�1@�B�����dV
'������7�=i�#)��z18�#���Frd����C����ZZ�u��*��=b��n+�D��=i3�q�{ms�`���sdz�I�t<��3�͝�^�ًmR�j�{g����jmtJ��t�z�tVř8w��"�V1�b8��lAe�{[p�mۨ�&Ì�o����g�P���m����-���(;iJ�^�1�ɂ��\/�������ю��t���ݞ�0+�=�j�n��nҭьv�wp\Av����D�u��u=ı,O�����ND�,K��{6��bX�'}��ND�,K߽�ND�,K�?G��-�f�f[����Kı=��i�~F9"X���z�9ı,O���m9ı,N�^��r%�bX���e�fe)n�.Rk5v��bX�'}��ND�,K��~�ND���DȞ�����r%�bX���]�"X�%����f[��[2K�32���r%�bX�w���r%�bX�����Kı>��ٴ�Kı;�x��r'�eL�b{���r�9s*� ������@�{��趹ı,O���m9ı,N�^=v��bX�'���6��bX�'����!�n�f���$c��m����q7B�um�181�vY$/<gKu�<s��9��9ı,O���m9ı,N�^=v��bX�'���6��bX�'}�z�9ı,O~���'��榵.k6��bX�'}��NB���'౯�Q��Ȗ'7��M�"X�%���z�9ı,O���m9ı,k�*�'�L�UH���Umpj�j}���iȖ%�bw���ӑ,K��;�fӑ,K��{�ND�,K��X��MQRD�D3E����Ibw���pI���͉ �'���pI�>�w��Kı>3�|a��\�3V幚�ND�,K��}�ND�,K���m9ı,O���m9ı,N�^��r%�bX���Y
~c�{$n��1�g�>xۧ�⃅T����<n9v{zY:vg���}�������%�b{����ӑ,K���ߦӑ,K���]�"X�%��w�ͧ"X�%��{}m��e�$��34k[ND�,K��~�ND�,K�׽v��bX�'���6��bX�'}���r%�bX��z�֜3,ԆYu���Kı;�{�iȖ%�b}��iȖ:Ey	詭�bg����Kı;�w�iȖ%�b~��Oֲ�fh�Y�֮ӑ,K��;�fӑ,K��o�iȖ%�b}�w�iȖ%�bw���ӑ,K���.BpѪkNjkR�iȖ%�bw�7��Kı>���Kı;�{�iȖ%�b}�w�iȖ%�g���~��ى{3گ<�Ը�^y���6�V%ۮL�Ä�ݤ,]���r�jx綵&�L�jq>�bX�'�뾻ND�,K�׽v��bX�'��}v��bX�'}�~�ND�,Kǽ�_\�j\��f�j�9ı,N�^��r%�bX�w]��r%�bX����l?�}"X�'�k��iȖ%�b~���?�	�5.K����Kı>���Kı;���r%�X�'��}v��bX�'}�z�9ı,O��BB]RSV���]�"X�-��xߦӑ,K����ӑ,K���]�"X�D<@���w9�ӑ,K����e�9l�).������Kı>���Kı;�{�iȖ%�b}�w�iȖ%�bw�7��Kı?t�����K���$�hѣzK���x-�|u����vD}����)�=	^yxՙ$�]j�9ı,N�^��r%�bX�w]��r%�bX����l?��DȖ%������r%�bX��ש�kZ�KsD�M�j�9ı,O����9�DȖ'����M�"X�%������r%�bX�����O���,O���.I8h�3FM]j���r%�bX������ND�,K�뾻ND�,K�׽v��bX�'��}v��bX�'�C^0��3	5��r\�WiȖ%�b}�w�iȖ%�bw���ӑ,K����ӑ,K��]D��?���Kı?���t�뙩�̸jY�5v��bX�'}�z�9ı,?������}ı,Ok���ND�,K�뾻ND�,Kcت�	���E;�n�{��~m���?Mb���z�#GO nT�������tZ![�\���F�6���}�ݱ�ۊ�c87k2����Uùx�ݦ�cvu�䮐��:�{N'۱h��W�R�u	�n[���;�85no$s�hWm]9�6�s��@��5�rFET�Kлp�;$�F�RQ��^,9�r*��z��H$��9�ϻ>J��
��$t�5/nڋ��-�:�ۊ��.q7��w{����{&�C���]�л��j���R��.��f1ǖ�k��*��zd2R<no�|}�}��ap�3R乚�O�%�b{����r%�bX���=v��bX�'��}v��bX�'}�z�9ı,O��BB]RSV���]�"X�%��{s�i���2&D�?{^��ND�,K�����ND�,K�뾻NDlK�������e�IufL�jj�9ı,O����9ı,N�^��r%�bX�w]��r%�`"{�����9ı,O{^?�.���.�0�˭]�"X�
X�����Kı>���Kı;�nz�9İ?�"�������@�o��_*��DD�$E)���Ȗ%�b}�w�iȖ%�bw����r%�bX�w]��r%�bX�����Kı:~��/�u30։u�����x^���Ȗֺۢëg���vܞ���bٕ�絣Ve6h�3NjkV�ӑ,K�ｹ��Kı>���Kı;�o�h�%�bX�g{��r%�bX��x�穔�Z�W&\��ND�,K�뾻NC�P�>X���t�'"X�׷ɴ�Kı;���iȖ%�bw����rؖ%��޻�����f\5,˚�ND�,K���6��bX�'���6��bX�'}��]�"X�%��u�]�"X�%���|L�Yp�3R�56��bX�b}��iȖ%�bw����r%�bX�w]��r%�b؝����Kı<~��		tR��fRk5v��bX�'}��]�"X�%��,{���O�X�%�����M�"X�%��u�]�"X�%�����ۻ���j�n�q�ut����ls�;v�z��=]�wݸ���ｮd���;���M]�"X�%��{�M�"X�%��{~�ND�,K�뾻ND�,K���ӑ,K��{���f���&�Y���Kı;�o�i�%�bX�g{��r%�bX���=v��bX�'���6��X�%����<k5��扐�35���Kı>��ٴ�Kı;�nz�9Ǯ�O� $#'�k��9����ӑ,K�����6��bX�'���KuM5LѓW5sY��K��dOr]�"X�%������r%�bX�����K��h���{鶸5P5_h��0OҦ ։��)��ND�,K��~�ND�,KｿM�"X�%��w�ͧ"X�%��xߦӑ,K��=I�)* ��s4�]O�6]x��m�ȹ�)W��d5�:�6����w�{Ѣ6�ri�O}܉bX�'}�z�9ı,O���m9ı,N���6��bX�'���6��bX�'�~��3�e�)��-���r%�bX�g{��r� ��,O��ND�,K�����Kı;�{�iȖ%�bx����5�̦�k6��bX�'}��]�"X�%��{�M�"X�12&D�����ӑ,K�����m9ı,O����yl�).�ə�M]�"X�(-��{�M�"X�%��k޻ND�,K��}�ND�,�`���?�Pbr�[��&sߧ.ӑ,K�����ֳN���	��jm9ı,N�^��r%�bXD��{�6�D�,K��۟�iȖ%�b}���iȖ%�b|w�ۿ[�kS!��te,�랇ml>�P:����4s!�כ��Y��5�I:鞅��d��5��ND�,K��}�ND�,K���ӑ,K���ߦ�9ı,N�^��r%�bX�3�}-�4h�3FM\��]�"X�%��{s�i�-�bX�w���r%�bX�����Kı>���O�2�D�?�r�al��ML��j�9ı,O����ӑ,K���]�"X��b}�w�iȖ%�bw����Kı<{�u��jfd�j���M�"X�,����]�"X�%������r%�bX���=v��bX6'���6��bX�'�~��L�Ys%3V���]�"X�%��u�]�"X�%��kǮӑ,K���ߦӑ,K���]�"X�%��j�CP�Ĉ �A
� sH�����'�ؑ"�BmZ@d҄��]>a	���\��5�߶=:BE�ȸ�2�:�D~SHH��E�� %JTp޶�K�N���+�N"m"@�"ET�`HE	6*���(��"�Fr��H EVVD� ������(�E�_�0dS|��	 A )-Dʤ�2�ȝꌐcCp�)���GR/��!wb��/1Ȅ �_�1 ��F	��*h�"E`H����awv����6?;��r�R�UU��p[F�[\  ���6݀�6�ˎ�W��gvŞ�l�#�lU@T�R1a�dո��� �.�(�n���q��p����x�[����E��.2��m�+F��.��WZŝ���69�ŝ�JKȭ�Urj��g�VC��ܝw0Q�r\�Z��+h.�i�d��&�V��{�@��Qg;l��k��.۶G�EL�v{b4�qZ+N�V�ji
a��+�^���[y1��:w��Y�h
)U�X��C(栬[�����+���÷n����:u���Y𴭖۵�5���[���6%����\j�sm�F���@a�(d��udkz#`8��;�=ttK��i�N��A��oF���@�v�l��x��kuJ�lZ5�Z���q�]�si�v�F:����v˪k�99��\��[2���<f����x����v^iZ!9^v��@WÖym��Y�kiv��]웑��%�z6���k[#
�`˄�MQ�*9����7n{3�IL�J2��;Z�-������ V�)�؃2��C��N���dzwc���׮�^�<q�@f�Y�Js����&N��:��TC���0 �j���9�^����lm���`L�.����(�ڕv�,2W����u@4���Uk$ vEl��ڶ(��H����[�\�J��e��
�yv��'*l�$�5�%�U�'��x(��%�[gP�X�v����fݸ�;u\�r�n����l�=;5Z�Vٍ��&3�����#]d��ML-�m��I6���4���(��(�*��|$�l�#�xx-��h��K\ݳ����6�Kg<��Ƿ#���xx�0�z�J��{=I�1���)b��fؓj�WA�ܴ
/7�٨�.ZxZ�zQ�[:�&�*�Nw����P �ل]���L՛��|"��k]�s��]��u�`W���3��|���ꄙV�p���; ��wm��3E��D13!�"�!����T� ��Tb!���WK�S�pS��hO��/�P^�!m?.�`M�q%l̑g���セa^Ʉ�J;ɪ�rb35iwk �֫��5�.w6��"�gm�㞞ܭ��m��N���c�^R{�Ŏ���5j-۳6R�;U�����=�ӟG[�.�Aݓ�rǁ�j��R��ٹۧh{hѵq	��t���Je]Q��͞���ywe���'i���u������v��øz�tg�3Ve�B(��������YN�u���Ҏ��ݗh�nq[��\[>v���p�ר���BB]��d̤�j�=ı,Oߵ��iȖ%�b}���iȖ%�bw�����'�2%�b~���v��bX��>�`�D��I������@�'���6��bX�'}�z�9ı,O����9ı,N�^=v���̉�,O{^?�Z�:.��&�Y���Kı=�����Kı>���Kı;�x��r%�bX�w���r%�bX����ƳXB��2jۚ�]�"@�@�woŵ�|9������-�D�,K�����Kı;�{�i������*)R(�RTIE�Ȗ%�bw����Kı>�w��Kı;�{�iȖ%�b}���iȖ%�b ww�����I��h.b�ר뎵�ݪ�7G�6F�a��v�;�ņ#�'���){;uv����{���7���{�{���ND�,K�׽v��bX�'���6�$�&D�,Ok���ND� j�_}⤢�HSQ$��mpj�K�׽v��柂�,��т�?%UP�r'"X�����Kı>��z�9ı,O���m9�2�D�?a�d��0����unf�ӑ,K���o�m9ı,N�^=v��bX�'���6��bX�'}�z�9ı,O~��		����S2��SiȖ%��"{����r%�bX����M�"X�%��k޻ND�,��~�ND�,Kߎ�e��[��Vd���ND�,K��~�ND�,K {�����%�b}���iȖ%�b{����Kı?{��w�Ze�uv���*]'Y�]��|Ľv{U�f���#�\��Ν#�n��ϷU^�ta=�~O������y�t׫����4���I��"j8�;�7䏾g�@���Z�Z��eDY2a�EQ`nέ�������8����ĥBi�R�;�٭�7kK3K�H�$�m�Z�Қ�ՠy�)�Z�U�\�E��q6Ŏ&]�v��=�{�Ir��?w������<5౑<1�� �Q�Re�=u;����v�{��[��':�{;�ٳ��!]��?w���tց���J��K�h�!AFX�e�Uڡfv魜�H����%ȴ��3}UT��N��J�����h7���֓�\���z�,����`fN-���J�*T�*�0��9T����y�tօ�S煮4 #�u�N��_��r�:��91c��MG��t��m�b��ei`n��X6�k�=�B �/m>�_�T�>��sI������\�ݸ��y3��T|�v�m�T�
j�TIG@�����;�4]�@�S@��㊩�HU"�&eTX̭/��M��Iݞ���O�.ɞ4ɗ�鵋�*�L��5L���Ł���ϛI��3��h�~Z���:<M��r,fV�wjv,d�Ň�i��}��}�O�#HQ�ck!�{�:�d�Ł�����������$���P'�J�Ԇ���ι!l�浙��a�NUUNt�F�M����c��WY��"�[+#�q�9�.�Y���kZ�fY�f���0�������j��ؚ^�Ev���ұ���e�y'v��:lP��GduD���v�����q����ps�햵dx�n�v$st�(��Z$�=��(snz�Y=� ii�9�0��a�V��f�.��0w����Sv���kY��mm�ba�[��r�v��rZ��#�2�ZH˻F�O(4����(�I#�����@�kK����'�m��d7�T��G��#��iA�#r-�������bG�ύ�eŠ~����+���Ge�^]*���!��gƁ�X���ߒ�� �ZX���R��%�m��n���ύ���<��h�d��*T�U"�D��X�V��i-��� ����c�@�>�c�6��33xc;.S���f-���RVC=������`["q7�2&�u����M�ڝ��I/�mvCw��`dh��O�L��[�njnIϻ���D>)�U�k"��k@��q�[�o���]���ADk�X)����=��4x�[)�{��<����I�L�G��ܪ�n~�{���3@�����e�9�ƣưrHh�M��_vl?�2��>����␱ �͐}���p��hꓷi�q���#ŵ�='g��{-K��J���[s`J�ͷ����M���3���L���v�UJ���B��,���_ɴ�A���g��z�q�3����I|��7��6ax&��-��Ɓ�ڴ���~N�	���I������ح,Y�R�j�]��������H��d4��3C�]��h.�R���uwu����h|���rV����hv��=]��\'��)�8�Ĵ@h��g��6�Ů/Gv2�L{��G'N��6�'��v�f�rVC@���:��������P�	Z�J˼��@�猿�bmD������x�3uV����r��g�2󗖖����@��yh{e4�%4/Jh�qP�@∫ĕ�b��䪫}��N��h�q��D��Lěm.&�S���X�05B�T�*�T*�����ZX5�I�}?x�	����߻��>�����_J��qw4��ćn����%pm�\g����X��(�FI��	0�1,p�<�)�u�k@���NW9����YӋ.��q7���p�:�V������ѱ`sr���i|�i��#G"~�"%]��ŠG3Ɓ��kOs�}C@r�Z��(e�ˤ*�@�UW*���E�}C@�և��W�8�~�/�bkF��E�yzS@�7�I4����tl��36�b���K!ZRN�%���,��Y��l�f�mșk�5#���
�^ώb�ֵ�1{[V۔�4H6����cU�'�f܆�n��D�I�o\�!7m���@����9�₯n�Ӳͩ�͆�p�n���Ƌ�\)���͵v(vK�����2�K�
��l΃I����ɺ���>Ή�ck���4�ݹx�tV�cS�K�ۨ6ll�e	���t��[k�=�������eu��y����Ɇ�2���tGQ�%�s��3�������.�.�ɡĆS�D�o�a5Ttd����lX�Q��m����|h�)�X���$��h����CsZ��4�mo���9I�\>�$Ƀ$��"��-�/����MܮU9�/�>����鎮��A�F+��[>�!�9r-�w���W8����BaVEx����.���h�Jh�*�/Jh��.�����N�\����`;��k��f��c��;�zd�^77﻽��?g�ìI7�^��@�U�yzS@��Z��`�x���Ru����~���J)j��X*"��`��a�@0��:�T����:h\�@���o��#��SU!]��Y��hG��:���T���h��@=��b�~Q�&��Hh��w+K3j6,>o�ۜ�����/R��U���^f-�w�z��r�������4�mh��
�ł�]�G"�Վ��V���쾠�"r��(�8��I8�!{�������v��Wm� ��Z��4�ՠw�w4o���I�M���@��������ȴ�6������BaVEx���J(��,n֖w6՘�R�ֶ��a��``t n�$�(6���'4a�� $�ե��O��Ε�͑� �$t|fЃ���~!���!��*�O� 3*Ҧ$�!&ך�&�v#�o{�H�b�A��y	��&ҘH�0��B!�`�H���ji��e��T �b�:Sb� ��h�
�J��C�N tQ8�����W�
!E�« ���t(�;8�6�S�7QȰ;�ZX��F�t�V��+2�+Bs��.9�@󘼴ϲ�����e0G�4b��'3@��FŁ�O��}�|t���9����������Π��&�C�6��zi4�:w�ܓӤ�^O�9���v4�pkr 1��&9"��=�|h�w4;���fg�>��@:����?(�XG$4�[��q#��ց:�E�~�q���RGe�}�,Y�"4������_z*�=����������&LjҰ�M(�mǢ��z�X��V	'L>��B	�)��	���znI��\x�1��0��Qhu��/��;���vc6l�{��"�Tv����68�Mr�m��"��)�q��#��qQ��6ݫ&�%̄T�%L�7�X��V;1�63kK���D�*&H����iX��W��mDɍ��9��?|���� ��(e�X�*����Vrc}63kK>i����{֬�����)Vo�L����䣻��`w=�Vs6Շ��$�S�q|��#s�Q5�rC@��V��m��_��1�M������$��w�y81!T@S ���� L��0�6"s�i1l��Snܕ��3�9ӴUӘ��gn#�㧮;68����n��ɷl���껣K�i��� �y�|�c�k���:׀��(�h�W)��M��6pi̪��j���;����g���mq�Bd�÷<��m��O/k9��ٞ���m3`C�hڗ�s�k���gV���9&��i륶��\�����3˱��{��w�0|��nz8�	Lmh�mv@�!v���4tF����晽��w���{����q�d��^(��hv�w�}׌�W��"�>��>��L��&" N�կ@�6��M>@g�ދ7����m��i�29�=WWxUҬ�1]��e�{<h;mh��uڒ�"��4�%�K��L�6�n7���3}�Vrcu����=_�]���ؙ#�-�NW9\��R_�:�C@��k@t;f�Oǐ�ђ`��<�Y�[N����>��s�>rmF�p��Q�]���x�I]�hv�w�}׌�>v��s��6� �E�Z�Ŗ��v�/@�����dȀGrT��?� �S��ܻ߯ۚ�;V�[S�I�Ll%��|�3@���i*�\�]v���O��}pNLx��(�Ru��ݴ��7�Е�r�ݓ�h��S���k��w��~��]���}�74�w4y��b�p&%$?'nh(뎴�v�����({e��ֶ�/;��a����j��d��5#�=�S@��w4���Us��}��Z�	�\Wv�!]a�4=�s@�s@���Z��o��$uq���t��/�.����9�sb��PД(��i`w7mX�v�e],.�]�]�hNR�����d4�7���M�����,��Z\$�Ye��7��'ݓ�~�6��Z��4���x��Q"�rDʙ�\�tY�X��'�Χ	V�#���eݥ��}���vI#�㉏q��:�nh��hz�W�Z���}��6�x%��7׵��vӗ�In-���o�UI��}�L��'�&�h�W�[}kOr���mh9��}�V:�f+��&Ac�ԏ@��Z��h��п�t��3DM�!.�`�5p��Ɨ���9����O�fb*�EL�Š~o�{���_�����Z�'��!땼�a��3R�!L���,Ν砼�qs����8�o#�^#�o9vl𠖑^��ͭ�����R��\�þ���L s(<X�s4y��@n�ց��f��^־rs�d����?5�i��;��;��{s@��qUv7#�G#Ǎ4��<�S@����>�}kBr�x��uqU�j7�Q4�4-���>�@�}U�������J��X7�Q� `N�:l�B�I�N�ҁv�{y��ڶ۱�ŢR���Lv��$�U�8���.1ɻc8�W9�;N�
Qo/4J\�ض�P�h���y��X$�=�ۉ{m]g�=�4��#����[�`���V����^�N�F���#��D��X��{/��nc��:����������V�8�ݬ�mZ����h�ֳQ�Oi.T'�!�-�{��ǿ�80u����j.s4�n{���gh�f�mN��Ϟ��2�g����M�I����ne�;��;�U�yl���s@��.<N&$ȓB�@�}V�岚����U�ܯUU�ڄ®�����Yv���{<h�{Zz��Yn-�qh*�]��]+�V`�J�Е\�UU���ՠ8\��;�U�yl��yz�Ŋ6�nf����;�U�yl���s@��P,��1A��?̚yq�6x�{=uً���;u.�>ѻ���eؾ}��҄����]�h[)�ym��=��Z�ջ$��#q�Ć��<�SzҌnדIM��vՁ�'}Ff́�҄q�r6�q�܆��s@��ִ�r��M��>�!�~��4a���M7SYs4o�6��A���w$����@��M�n�m�f'�D�c�RMTX�6ɴ�ɴ�}�>:}�mht���{�TWK1ave�qr�9�0��îS
����Ru��r�A����N-8��Ǒ4H��c���}>4-���>�@��^����0u�<i�LJ��?6�����UR���ZRz���h{n�`�ǎ6�nf���ܓ������Ȕ��"T�"�*��ǲ�v��
�!��ikV�/�m$��׋3~�`gp"��6��hL�n-�uz��h[w4Ԕ�N�vG!�5<HnM������M���4�k>���+�@��^�?g:� 1�a�O�mD�ݪC�j���i9g�^�h7jGc���%���tU�GH��ƛr�빠^����3g�&�K���Ł��<��H��q�Z���Y���z��z�{��@������)#�Cn�լV
�����@i�zo��\�*���M�8d4}�#Ǖ5d#�@��h[���+K�Lm!$0nD��$�*nP��I��^�l��'�N4�&$�ym��/RS@��^�m�������\'��(������o�G?Wiv���b�����^t�ǋŶe�u�b�.�]�]�~8d4�]��g���s�	��b�
��-
���0�?�R��	&C@o�k@}f3}\�q d�]̵��̻�V���I��빠^���U��}����D�`�����s�G?V�2O��<�i�?}�>,Q��QR�R"��QDL��/RS@��z�S@��怷��2G��:n
���c߾��N@G2TaYI�S퐋 ����Y�Ke4�2"���	c��! &�B1B���M
.�b�CL�U� �ڜ>�~OBsZo�N�	��|#���WK���$M�44I'��(�["�jHA�~(<a�!�@/�w�?O��dYh�lm�n� 6�am-�8lޡm�`8��l}e��Q�r\i��H�R�n�fg-�vE�{�)�\�Ҫ��%c�t�-�$��G\�ڠ�q3\��M�����.�z8��ulI���Kg�S�Pm�%����җD��v�Ò�莈�g�˃4�1"+&
Bj ��U[U��ܹQ%E8�pvw+<fa;`j5F�ƹ�c,�R�۵8���;W/��e�G4r`��.d�l�諶`�h�؀�O�vv]����[Rc�&�U��b�`�
�헊�x�6�S�z���t�kn��"K���d˯`g���tc[<�<J�l��\A=�h�[���E��T4��"�\��N�ud �O\�+�j�I�ێ.'nye!�<-����Ѽ훗�Y�91xzw����Ջ{�(:�3��G�^H!���l1[��[���m��[](mY���&)�:2�U;�Y�ΐ4�u�Nc�gG��-��xHv�ۯfxv��x m�[x���ir�;=�����T��g e�G7Q֞8�2�3f�09W�ٔ����݌�uEʥUT�m���d%�L�u<\`s�4+Ue��7SUʜ�h�6Ŏ�v�۔�M�k����U��XJ)#�F�e�iykj��� r�XlV�6�OLX:h�z��N+[R��ڠ*�v\%��2t��ݷcA2I,UJ�!(s�[����n�rP��v�#rmܱ��SK�+�q"q�.��c����+�9�=R�Dm��t�ۜ���i�UV�L�D�����8�0+�T�^Ȼ��wgZ�k���%Z&4��l���1�Z����rn��x&��#�i;gψ�L;<5�j�F�����L���*��=���%��\g=��nʝ'�[N��6\��T�R6�^v���m��a }�k�KT�:W1ۇ��Gj瀫� �l���Nr�d��Y*�W�6j�Η�sR˩s5x�At��6�( |�����/���(W�Tb"Ĉ���g®��8U{s2��<g����A�NBd�z�nZr��%zr�#
##��SVƼ�㓈��6N��Ͷ��:;r���k��S�6��]��1K�^g ]c�x���ix�Gg��s�l�FY�q�N�7:iwM�h=K�0e���ɺ��ͮ��z����͙��.�q��I�-G4+����)�s�����N�]ضۛ6ܻg�W��V9E&�v�������{�����,����N���2p^���q7�\�p�{vM�hWZqŝj����1S(�h�2;�6��Ł��k���_Xzx�u�.���b�WXf�z�ՠ[�s@�IM���߳1#՝*XZ��һ0V+�Z�mh��h^�@�ڴ���0J0y��V����qG��r���ʪ���رB�is��/0�4�]��I�/�H�ր��f�9NW�>w;�n݇r[����8�Ǣ�3�{]��0^
��]�۱�s!�����[��֧q2�V�������Z}{Z�1���W�}~zw��ȁ4
$ܑh��|Mq&�k��K��gj;c��`n�k}�H��d�.����8��]�hL>ZW��-v�޻���^65<X�M���@��z�ՠ[�sBr�sTZ�C.�+�XZ��,����ց��r��G>����@i���|��߂��V���R
�u�\m��xӇ�����S(��#��77�������,Wx�ޞ��^&��]��V���܆	F#�Bnf�y�k@i�ހݶ����$6Ŋ+K��Yy���r��mi|�r��
� �!�!��!H:H��H@�� �.N�C�մN��Ձ����a��6J�SSS*�3Sa���BMϽu�$sk@m�4%r��~�O^�߱z��2��4
&���o]��)�Uz��)�^�G�����"Y��x�����A���Ռh��c���!m!YrB��o����0������ ��ƁU��l�����G6�	�We����Yt��4��g)"I��$sk@m�7�H}�,�Eyk�a�^e�L���^֞�s����(���|S���+�y"���o]��)�U�C̿��nRT����`w6����UJ�	���S@��z�S@���ߟ�8�ߝ@آ�o8m�u,����ݿ签ݶ��ަ�����^�[�-�XKv�;��0�Q��x�����? �d4
���qDc�,Y1Ǡ[e4����3@�}w�ʮr�Uv7�U�3^Z���4	���M���Us�ʤ��^�$�h�}x,2��YVbĮ�'�a�5��mhJ��.z{����x�?��r&�'���W*����sk@m�4U\9(% ��,����'�Ժfe��Xک����s�֎�i�Br�:,-�nz��h�'����!�{9ŵ�`��7v�2�Lvs�l֋m�wV�O�s�y6������˄z�����Uc#��*>]�[��"Si׎5�&.�:�=���d�$�3mm8ŗm���Vޫ�����mq.66��qg3p�l���a�Dե����z۷\�9椺W]���lu=�F0��������i�K:vH��l�3:�1�n9�Z��b�'e�=���NCX�OIu��j	)#����u빠[c?����^��,-JJ�]�+�-�]��)�r�^�k�h{fS��xchM��/YM���Tw"�$sk@�z#�Z\�bE���h>���$Gr-G6�<����ؾqDc�G�<Cq���@��k@}x���z�\���Kn���n::wf�{y�����]�w]aSC�;vF�v;�f7�q:���6!&?�o���߻@}x���~��܋@�&%���T�)*(��V�֗i1�%�)IbeS��<�j�-빠[�x��X�U�+��4��@}�֞�W9w�Onh�O�@�r�4Ġ,qH9�yڴz�h���U��q��c�]W�X��h��h���G6�����ՠyC�Q��-�}eB��2)����[���'=ps�<��(=u�z"y1(ƈ��Л��^��W��/;V�o]���J�C_�bC/30�}w��U\�H��Z�mh���ʫ��X��x$�z�lX����mJE�BI	&�S�k��+�����d��\,F�f���F��X^Z��^-Ur��R��ՠG3�@��z�j�<��"x�!s4�S@��z�j�-빡���'��6L��2����O�tux�	�}1n���wc@�{8�}��{�|�\���&	��>__��yڴz�h�����h+�A&� �z�v/W�I�2g�J����X{�_4�A����e�< ���@����/YM����ՠy��0ʣ(���34�<�&�J~����>���`nN�Xko��mB���'us�Vw+a1�bC�^�z�j�/�w4ͭ,�I��5z�*4I5J;]�E��u��6R�q:F3&s[gDsi�uf���f~͑n-n1c�7����?���@u�h���"뗠>�S��/#m���@����/YM�z��o�~��H���AH�,C�E������*���/;V�}빠[�x��X��Ȕ�U�W�^v���kBs�ʥ�h�Ae���`��3	#�/;V�}빠^��^�z��{�ߝ�m��[�&ܻ6�1Qm���je�^ȩI��㊶y��s3K��"㫒6C��8��t �onr$�����{ǋ��/\��{r�ر֝˫t�KC��lic�7[�p�f�l�-�N��n��<gp�m��%�w=;3l�6m��;m����|�啐��4#ˍ�^�k�:�aZ:�E���K�]V�,<��3�5�! �jh�������y�u���\��&���.2M��!D%�s+����C���M���z��s��/'\f
�w��G��>�f���W9�~Aȴ�2�@,B��E+@�+@}x���z�����ʪ�q!�,P�Z\�bE���h9/@}�֞i��ʹ�~��Z�>���`��fiL'�(�ǈn=�h���/YM����;� $���%Z���UU{�UU��}_�=��m���r��C"�����G��B�O��q�[rKqF�f��ϞN�P��3���8���[f�z�������@�n�o�x�X��7�p�*�^���1g��LD�(T����~�~��|���^3}\�U$6AeҲ``�Z�1f-;�hm�i+�G2�$X��̐�LJ����&j,<�m6��{�V��{<h�k@n�ZP
$��Ĝ��)�{zS@�ִ��ց��Ju"*_�.쥂���'�M�/<�v��.9�{8�8��y�h݉�}��vOS��O蘐�䇠u��Ɓk�h��s@�e4��U��c�xc�ۆ�z�h��s@�e4=}V���g��D��"A$m�����=��恛����>b���`�ĵ	�q5�A`O�S�@!�U����!�١�$��_�$KA��q�4K\��an�S�d�5 � Dx���N<��9k��a��4��0�"Ă�"8"o3N��e�t�b� ��f���`�4p�+ ����p��)ݖ�f4)nJa��g�@���)�8�YO�~Qu>P:���������|!��D� ��D�.?�����8�~���y�$IE���U�V*�RW��92ﯭho��W�s�h}H���7�r(М4=}V���h����:�3@�*BjR��X]�u��-��7&�r�V�R�vKGDs��-����q؍�M�y AbjE��/�O��͵`f�i��IvC6}�XOL��M<M�LI�@�޻�[)�y��z�h�2��!G�&�'3@��3@��q�N%�2�sk}I�+�ȕ�H�H��,8�j;�~,�W��͵a�ڎ47�_!)I5ƚ�ﾭ��}���5�Qa�#��e4�^�u�~��9��~��� ������~������;�ęM�6�+v��i0�<�`�^9Κ�M�UpV�m��?��v��YM�zS@����n��őՊ�Ŕ��hu�6W)#���h{�s�#�H�<5��<��'޳�@����=�S@������`�Z�Y�����M͆��\��=�S@���h/O�ز�O�`�;�j�������p�������O¿(|bT�C&��7Q�,�!���Y�$-��\�3�<,;���༵�zS��r�3g*O+�\,o1�S���W����S	7Eٷ�,���H��xE�n,l�ڎZ��l�o��*��)n��c�
+�5K�Z�wiP�Ϣ�d��Y�����@�����ڢ4�L��˻-7bu��>�d�y��\"'j����x�	�\����Jy祁� D��Ɋ6J�II�g��y��?tp}��㑫�t�/c�d��t��ې�/ˬ(�Bˢ��%yP	�g���ذ;�Z|�|��o�X��M�"R�ܐ�<��4m��<����n�Wu�&��,G4m�h����r�UI7&ց�^C@�牲8��#i�����w4�w4=�M�e4p}`����D����ݵ`y��o�� �z�Xͭ,����3��Ӻ{V�j�cp�(ݟUu����=���q�=���\:˗��8wf"�N�e4m��=�)߳?�33����>�]]���R���/��]�ҘD�E�A�N���i�M�$�Jh���X����;�`x�?T�eƞ&�'�p�=�)�w[���\��%�r-�d4��eeաe�Wi+�4%{��W.O{���x�>�S@�����=_�i~��nHh]�@��M���;���nrJ����loW:�Q�j�Ugr��y:��+���{'gmۛMv�{������*�瘎�D��p���������i�I4� 7�~Zw�}�90��D1I�ץ6W*�ćِ���󾵳�ʪ�;�.{-V*�V�+�4��4�뻕yDO肔����!�6����3Ϣ���_�
��fJ1ȓp�:��@���@�Қ{e4)E7�&��8�k�	U\q�? �2]���UT���껴j��+f��޼m�J��<�V9˳m�c�k;��H����<u���E��>4��h_U�{_U�y�R�QR�3TXݭ/�4���\���yh}�o�#�!z����+��/������:���ץ,Ff�UU3U0�TLUE��M'�MO��}���,ܭ,-5�!�4�f�B0I��&"xB
.��@6�&Ǚ����w��ra����1I���h߲�w��/���Z�y��3$�6�''�Օ�	<��E�j�4bsӸ�g;d��\�+���1��(,c�	�x�ύ��h_U�u��{�x�5V"LI�@��Z��Z[)�w�S@��Y`AbjI�@���@�x�=\�9�W.�x�'��Z�Ӎ^,��<O$O�hl��ץ4�����sZ{2�Eb��/
*�%y����f��q̑~(��o�k��8����um�%5&HLu�Ӈ2�c�ݣv�wu:;�tOe�Ů�g��etdF��P��

�����*�����6#���эg�ـRC�q��\ñ@㴆���:)1�+��g�!ӛ<�Ж�0`ޥ�w��a�6���%e�
��|⺱s��L�m�7*a�Ǌ�@���*�c�a1����x�u]��v�k�Xo&M�-u����ڥ3-/��v�_(A����&�UT��Za�ⱱ����O����5�p�x$V��,ǲ�˴%e�f���R��BW+�	C@�7��eX,�T���Š4��g?���O{k@��x�>v���B��q�&,��$������h����v����\nPXǐ$�h����v����O������_���<�0N�ڴ
�W�w[��[Қ��U�c�I)ѥ8ѝ���ˢ^ۢH�$vX�`�{p8��%�]�<v�֕�V�8J���߇�]��{Z}�J��;.E�|��v/�*��b�l��W��KM&;�\ύ�r-��{䏻2�Ee�Wf*)ZB��vd4����)(���[�ۚ��ՙG��m��ػ���"n^�ߛ���p���4��̉L`�k�ԋ@�����s@��M�������#O���,��=��ހ��#��qՈ�ɨݐ�]̳p<����̉��q�$x��#�����~x��}k�~@�Z�RD�\�"Պ�y@Nf�m� 󟼴]�z{^����8nR�/
,�Ĭ�v[�ܓ������c ���( H� ��A`�BՁR#]M4�����M*Mv����;����R6Ŗb�Ԓ)�B�^���j���ia�k�s�_��#G����j%R=��s@��M������hv*6��ƚ�X�!l�rh�BE�j�+v��ps�g��'#l��zݺ,����_l���}V�Wuz{n����fF�BLnHh��o���r�Wg���?{k@<f��w�I�F�<MH���=��s@��M����lW$r �$A�UM�ͤҍ�{���z�X�͋
1����oğ֕��N>�s�>_ÿ�,i������e4k�
���;�w4=ƪX��BRd8�ٛ	k�t�n+�����b��t���7�8:
�Ìg�2LOD�����}V�W�w�w���+�ʯ�'^C@p�]تe�q�E"�*���;�w4��h��h/OձPi���D�@�m���^i*�UĻ-ŠE�/@���26cd@&��� ��h��h{k�<��h[^���##hI��M��ZW��<��h�f�q�x���Ni�!B0a�@d��FHq��,�KYQ�!�(�G�]
��A:8�g��WF���ة �07S���≼΀@��4�A)D4��D�X�o� ��I�����!�)����6�9���k�Sڹ�*V)�W� L��ç�~~H�t	�]>@�E�(���B��*��}����>��I�:=�?_���l�`���v�ڶ�6��� �W-X̙���^�q��A�6 �^��jV3�ٹ݂n���Y����"�<��i4����n�ȶt̺����m#�7����ۢ�<�4ۃd���EWV���7e&�ds�Xؠ"x�9���ͺ��Q���"����R�S�R�m���ԙէ���g��D�v��T[�(����h~q�*��AE�oF��6��=4��iBshA5�:�n�p�[\p��h�T��xУ����j�5+��A\( 6d�n^2F�@����`�n��������)v+�ȸ9���`-E�ܝ���2Ӷg��»���
��Gsd��ͷktm�[���1���(m>��հ%q%@�s���˚t3�u�c�6�'L<p���rkE��ns�+��ɲ��;n���V�E�^\5�ܵ�u��gm��b8�	4��F��veڥy�Tp6�9iV79���q�NY.��듷
q;�s�U:2]J�.�q��{~���n�"/����ӒM�����ѯV�I�]�JQ��I�'�q<�v��6L�����@��ؼoK*�US�9�`�:KvM�W�5&�V��+ʭN�P���X��� �n@.�ˬ�	V�PVz^V���RJ�o0[@�l�mq�m���R�ւ�Ӛ�H"�j8%� �Mu���/[�Yɴ�>����z��*�JA���Rm��Rqg {6��c�/j6��pu���Y�6���6�Z��%�&�r�ɭk.�ĭ�gml��l�*���=��۩V�c�&E\�Ә���T*K5���7d���5��w.�b3��V4cM��/v������JF��qYm�>KRm\m�*�i25\�/U+�@^'��d��{,��0ή�6����m��%LT�/^�K�Ym�/ ''@,R����&[zdv�ge�ۢϲOo?ރ�Y4s�
v�ل�ju�)�X�ytYē�mM%�ե���5(�@?*� ئ�Pa^0��1AH�]�D(~qD:��ҝ D������j ����]�ؽ�uM�a��<���`zlZ���'��9N�q���ΎŭG)�.%^嵊T�8�9GT8�7�o�Y��z*H��;[lV���j�֏=��i�ƛ��')�7n�ssld0��P�u�nG�;�����m;.��m;s�nl;v&yP�O�u���p��M�l�e�:: �����"���U�7K���D���QB���2Q_�k�1��O���:�����a�H]GE�H�ۋ��]�0�P5�\�n�6�����}6z1	����MH���w���<��h�f������XG��FG�@�۹�[њ{}k@i���+���]���ؕZ�X��J"iX}���3'6,�$�Q���I6����WW��X^bX
��;��ZO��ͽ�UR��4ψ�}@'$R-���ٞ���_���%s��v��>CeJV�e�y�N�w;\�fNhثw="��+�뎻ѲE�L�F����@i����R=�n�}��s�
���=�)�;!�M�).hܓ�w]��q�tU�4um���t]N�,Fo����ڿ�m%{����J�4�crC@�ߖ�Wuz����e4
�R9	A�ҵ��')Kn^���k@<f���Z�=��`�`"F�Yr=�n�oJhl��U����������e���e�^,J��mё`����ɶy0�,�x�$Ki��G�9��)�u�f����~@��h8nR���J���+�@��3g*��"n^��ύ�e7�H����}@'"��w�`f�iga����Z�I��_���ύ�JblTi��R=�Jh���ץ4
�W�y^q�"vI*��������$�{��~(��}�h�u,+Veݪ,3�k�"��q��S�����NC��<Y�lyqf(�1!�I�Jh^�@�Қ�)�Um�2A�9Ю��}w��ʤ�C@��4zS@�lV
F$x���#�-�Mޔ�;�j�*�^�s��ƋJ�3�.�����qH�]�����nM���AP�X"0� ��T�cA J~O�r�߼��;��J���+�K^/mzW��=�)�[Қ�K�(���q��ErѮe�#čcv������^�ۆ�z�Z�%ݱ�si獙�SZW��=�)�[Қ��4)��Pi���mH�oJo�$}��{女U��+�a�udcłk�4������r�(���8���՘��#X��$��u�4
�W�u�Mޔ�*�������@��z^��-�M ��hM�E�E��N��o�5$��ܤ����/��Δ��"'�힪p��p=0V͹5ؒ�K2mH�6�n�7Ka)ӯNC�Ә�v����97YCV9�+m����:m�����;q"m6x��s�㧲G�(��F-�gŸ�:����^���.\�8�Eڸ�(9P�u���of�{��8x�aĞ;�6�i{r�v��ά�2H��kt��m%�Kq�3Ɯ����?�����>�X`f�3j��&�Y��8�F�ͭ�Vvk��s��r��s�4�#�H�$��G���?�ޔ���\�Uj�]�*�T�+Ī�id����>�ύ ��h^�@��fĉ7)]^Z�ay�`+�@M���zS@��Z�������1�RM���zS@��Z����f��)]��Z�j�v�/@�Қ����f�U����0��w�=�g�z�������g���q�Ή-�\��yS;�$4l����[���㰝����|h^�@��_� �f���p�T�T$����3sj�7�&�I�?��'����h��h6�e�c0rO�NM�mz^���ľ�|h��4��bR #X��I�ץ4}}V�u�4���c�Y$����4W�^���~�O �w�=�JhZ��A��G��&9$͛��"����[C���t3�25��g<��F2C��LOk�'#��f���נu�O�fx��_���
<o�Lx��<�I�x���zS@�{��^�@�zSƨ$�MB7z^��=^�sr��!��I��G� |hC54���jn��g=V�g����q�����@���h�z� ��h��ބN=�����U,��-R�k���Y�x���zS@�{��v~l^w~;aܭ�SѺ�x�n��9-���Nt���[g���sa�	ژ�ݞ���94���Jh�z� ��h�+��3QI#�:����˯�@/��x����w44�I�GJ���]�_^i�%�엠8���lq�L"���C�����c=�;�ZXJz��l�$���� J��Q-�,!B�Iծffy�y}���F�H�X�Cq�h��́�����w6lf֖�i�����~�h���f&����D����Y�.�ۤŗ)�;�kD3��w}�����`SMB7~����������/YM��@�S N�lh���z����S@�{k�/[��ymz�y��J��Wyz��h��ޒ��M��_��˺��i3�M��x��������w��W8��7�a�018DRH���h�z���E�����Pۑz�$�ۆ�c���߮�&�$d�V����}׾�?d�M�W�6�[^a���p�vyv�cI�:P��R�l�r!r�˴��i޺ܵ���T�
��U���/J�NRg2nLM�gd*�Ygm�wUK�s=��:�����`1�� Q�׫2-�CV$aٺQ�݀.��y�6��VʨԦxC��G���H-N�g���	��.��� ��jkZ���W4\�4h�4K��EA绽�����?�?��E��]�T']���}�2s��<��2sɈ�8�Y4����vyI��	��=_���@�e�@�{k�/[��^�l�����)����\4������ޯ@:���R(	8��s��@�n�����/Yp�=��1<j���d$qǡ�g8���h]r�׎�	K�엠|�?�ɍ4`�Bs4W�^�zˆ��������
^m/a�#�I�!8�4wn]��E� P;<����u�ݽ���8M��Ǳ����,wݤㄅ�����_�����w=��@<^{�@�]ն�i�9����7$�������Q�v�iZm��srՁ̜ذ76��Qoĳw�T�Y���G&ց��ڴ�\4���Ƹ���m�b���w���/Yp�<W��:۹�[�ُ"���S�hl�h+��m��;��h�B��� �v%h|�1�/k��R;,g k�Ä�{�0���ە�ey-p2�Wo�����������������^q��W16AƤz�w5bG�������^��y� �Zi�ؓ��yӛ�֢ͦ���δ�H�m9s2Ax>��	�@5C���u��U�`�@��!$��pHG����2���|P�yC��8������H	�'�HJ�� �B��sBl� ���qbB�����L�C�����~8~"o�7� 2&����"��d�5�������s��' gM~�$��q�5^l�6�dV$a! �Ѱ,(�	#i@�WlƺM�*D�1
D��#vk�BR�����"���)�N)O�MS�!�>��#�o�;�I����O�pD��L�`�A��@������;�GD�C�3?RC��"�"������$�|�~vl!V4eHQ�Ft�N�'�|/�T�:��9�4�O�~)TND ��u�� Gmꁠ?ϟ�L^�D����v_� ���>�^���Te�T�,�š9�(��4�r����'+��/�@����$m5��1��h.��m������ˆ���e+�N{sջ-��h6�t�n�3��Dd�k[6{=�R�n\t��Eܶ�tM?l|���?v�ց޼tO�>M��'J� 4ӂ��I��<��h�\4Ff́�ݵ~m��A�o��*d�D��c�h�>�@<�@�۹�yϪ�iF�5H��r5	&�u�wvח ;������?C���P� #$�IH"b`H�Z�A1�����2(�2>7ZE�, ��P�|?���=��4�����1�A�������}V��e�@<�@����8�v�695�n��<�����|=�,7b�|&<����>x�;�å��
w��qh��F�~}y? �k@��{3y�k&�n-�ˆ����ă�}V{޵`s'6/ͤۈ23|MUL�&� Na����=��hs��.wEbN$���HܓC�ʥ�'��>v��;׎� �޼��[u �l�GNf��>�@���ڰ;���$����G������ݟJu.H�[ɸWvڴ�#�b���]���6��tU�,�0v7�4��/�
�snW8��"Ocy����cMm��6Lmڃe�Ngv���Mi�9�^�Cv3F���ng�2b鵆�������.b(��X7�kM��˷�d�x�ˑu�ެ�b��m�N�ܛ;���5�0P�Pp��n^�6�M�U�s��W���Յ�u�W�+�o�\��~� ��r5ж��6��'79�I���:�3X�;��u-��;���]��sG�m��~_��u���hs���o� ��jL4uz��h��l�o��#���lk�,cl��H�	$��;���%r�)&J4�r��q��ʘ�$�'3@�_U�[e�@�^�@���ε��Q�
,15qh�p�<W��-�s@�_U�{���l�=�t�;f�	�����v�B*���Y����%�t��wD�Z�Eݎnbi70�<W��-�s@�_U�[e�@��\�ȃ��ȣ��۹��'�D0Q�j*C���}����F��>��=:VK���e�'3�/;��-��x�W�[n���.<l�EI�H�l�h+��۹�yϪ�>W>>���RL<�o�@����}V�m��s��B�ڣ/2�����_����J�U��vQxoP�u<q*��◈|r�sdjG�}�ۚz���.��z�q�<���&�9�z���.��z��m�H���f(�����l�h+���?��B�i��6���Ձܝ�X��� X�14��h+��۹�w���-��^�E$��Ȳ�/@m�����q~I������;ӕ�5�X��4�,q����odJe����8�zn����&�4�7����hC������_U�[e�@�{��۹�{���Ȁ� ��h�ʴ���@o�k@���R�� �˫S6�9y���z�w4}}V�k�@�����T,cl��8�{mX��Ł�8�,!4����M�g�O��M{f䟏9�ɗ%*V+��?}}k@�$�Q~��/@o�s@��1��H�X�&��Q��K��7Ŕ�<�:{mnp%O@�c�NG�{S]��
,14�qx�;�-��W�[�s@���h��� X�14�ȴ�w�7׵�~��ր����U�$6�@�<#����������_U��In��>]r��ZlČ2�`'3@���h�p�<^�z��h���<�	"	�Z�\4��`n�ڰ9�͋�7hi�֦��v�˭�v�9���mL�tVƃMsJ�2O<�[Oc���;�%ڸ˹M�ɜ���{w��( �m��3Y]��q�;��-s2;��:��d-�6��,e�{v��n��mX����Y��X9x�ɝ��<h���m��;3p�;V!�gl�����]�N��G��콠��jn�����]n��k3��͞ģ���5�ܜL9��������w=���� ?}��\˭f�d��[%�͛�1�SmV���von�u��n83O�ŧc<��rC�N)&����۹�y��l�h��~�c_!ci�8��>��4=}V�m���W�yCq�cˉ��19����@��F����u��$�k@��w�T�ꅊ�M(�Z�\4�^�m�����@�VȠ��&�s��@m��ﯭh�th��Uq|�1��Wm�n���FC��Trtd�Z]�.�Xk��p8��|�S��f��u[�Y�`�M���ִ�:'9��\��W���j�8��m�����>�����Ip��H��� A-h�T�ʥ��衺���E�g���-�s@�A�<�H�F)�m� �޳@����_U�LW4��N)&�f�m�����@�ˆ�����I�H��-�s@���h�p�=�h��J��C�~D�A#"���j�BcՉ�2Ì�n�q�G����K�ܦ�s6�[�9�3�� �w�[e�@<�٠[n�綽��<�5�Q��m� ��f�m�����@�VȠ��1���"�9�ڰ7wmY	4�]Bm�Bi�Z8I6�ƚ\m�/'y�V���͸9D�S&$����-�s@���h�p�=�h\u�$M�b�	��=��Z�\4�m���ho���߇|X���V��3��/^9amԖݶr796��x���nҝ�����{<��L$ƤZ�\4�m���h��� �b�؞\`8D�a�{l�$[.�ﯪ�-��{��ccTi'��G&�m�����O���@<�٠yA��yq1&���h��m(̭�X��Ȱwv�!&�R�4����j��tٹqR�S
 ��f�@�ˆ�y�@����_U�{r����v�玣i9y��n��*�Y6���70-�ն���l9#�ȕ8���-ƀy�@����_U�[e�@�]��!L��ƛ�@����3=�~Z�%��ؑ�쬘f%�V��X0�f��Y�[e�@/�f�m��~t]��/,3��Bs�L���\�����q� �Ruv��2����Z_uހ�9\�*I>���>(��Q`|�i4�o�6�M6��ɢ���DU�0DU��EW��A_�(�*�𢠿� F
�* �D`�E*
� �D*�P �D ��H*U �EB
�E�� �E��F
�*�� *
���H("��"�"",��
�
�F"���
�H* *��A��*��(��� *� �B"�
�`�AH* ��DH*
�D�����������H 
B�*�
������
�� �A *b�@ *���
�b* �@��@��A��"�`*E �AQ��AP��@`�D *H
���2( �H*"�DP�����DU�uEW�DU� ��EW��A_�QU�DU�uEW�A_�QU~QU�1AY&SY�X�]�ـpP��3'� an�      �   �    ��  �� x  |� P� �A@���    (�  �!B"
@     $�   " �   # � �c 
篩sof�&�eɥ��-�o �^���so^�z=u���Ҹ@3�X��[����o��U}��W�}� {�L��eͫ�{y4z�6��� ,t�O6���}�}���� �   <  ( 

 RVX S�'��r�[Ө��ʽ� >�gԹ�֞���W�[�:ˀ6�w7R��v�i嗶����� ��+�U;�W�qizr�N�� ��m���U��R㻥��|ܫ��}@PH 
AD� ���Z��{ݧ���:R�\���г��nR���R�14����J}�K�R���)JZe( ,����YJ
X )JR���R��vR�R�hR�=��)e��u�(���(��R� \r�J @�E� �JR��r�R�f�M������� ���Z�9k��w����mR�@ҽ����� Mũ�ۥ^x t�W���e{�u{{���y{����� >�Jͩ����n����m7�> 
U( P TX�Ѣ��_Vێ�^��v�g��{{�[�Z{� {�����R�^Yy4����um��g����ｹo7.� ��ޭ�o�ξ�ܠ
M*;�r�9��qܯ'.OU��.�������^,�W6�V㺕x   ���m��H@A�����ʛʥ)P  "x�T�5L�Fa1��R��IH  ����T�Pd21DPLR�@F#LJ��?/����?���>7Qo���I%
"��_� Ur 
��� *�� ��P EV*�������P���`ɦ5���?�pdaF� D0X`!�pE���O�)񙿣�Ϯ\�"a8�9q!�2�
�A�\00j;��CHD 96e!!P���eqE�n�Sa	7����bH7iM����b�%t��H�ha���B���0���)�D(K�Is�,�
1h���\�e0B�x�eaD)\9p�{���kgS����}'�h���!bB6$��9�0��lp�_�4�SN	�!��0b��� "��HI0r������J�V�dR!�0�t��Ϗ�ѡ�FF!#�J��@��̃B& ��r�"cB^�e.�V;��֛�BL`�p�[���F�:2|�%+�\d6GaW
� �� ՌZr�c���tL���B�! `s n6C�M���ʄ)�,h`X%d�7�/��ώ��Gd����d	P��`L)��N����MF	.Č�dFI���N�@�d�M:�~N
�#3��}F�2vB$Z1	#  �$�2��L1��0!! ��B�@(hv'���|!��Z�
8>y��b�I(a�pٛB�պi$�t�8�B��vf����+n�#��)��e���a!H�H��pTs!$J�
��I	��#���w
�CSDƀ�lhĀ9H��T0�SΎo��$)3������*B��\1z��b�bW��C��&w�@� �R�S��cr��H\L�B����q�Hg&ΪcG��0 A�J�$B�E�A�Aq�C;)�@����\$`T��eL�����۔�BW �b�̑,\	���e�h�
d!P��Ȅ�� d�p@��$~vMo�>�J`������H���L�&�S��/^Hta\�AR�XD
e���ii�*��	&�˃&8p��Wi!~�vfdɰ�A�MZf�f"}~s�dː�3p?,g�B�3:�՟gI2$�>yV�	74��X#��W�㋩>D��Y���a�"� �U��;���`X�$"%"�	h�	�n���G)$�ߤ�m�L�
r��l��Y�Hl�R; IC5��� U��R���`�0��\I�����d�Әh} ��
"a!T�@��q�l�R�B�,��"H�1&��D�2pÔ�Wm%~��!G�.\�!�!��!:���h�":�����C̌
�2e��~/Đ)���,��c ��1�sM$@��Bp�t
`ɠ ���{s������ @O��-@�L56g�����u3��Ӻ���X� �"��"S���(V�D(�"�		"Ҝ��B��6�b�@ d�rF�}u�T� � �*A�$ v�ۈ�.%1�̛�3Xϋ���� iupَG;ܲ�vj= Ә�Lh4��|��$1���J��: ϡd�X��%���#�Se��$�a``209c�����X����1�Q��X@�\�|�;ӧ���1Z2EH��!q$K�LJa��.pk_����F}p8�d�*P �S0��]kn��&rg6J�D2�{ٰ�e������ù�ݔ�,Í��wX���R��nf���(�9u�%��1�g@l�>&!)y%#���-X��� Ȧ��iȑ�/�W(�)m9�4���w�Y�\)����9���C��.1�B��LL��>���Wa�đ0.$XBG[#L�z5��6:H5�#	P��H�p1(c�p�U��ϱ�"A�E�Pљ4��u�SI���i�b, �H	HDp0
�"- > "X%D>e���}0�9�֍��!�f��5����%�����!�A*��S�P�C��j�ӻ�sf��0a�0C� ��e�����\e�mK��0B����0/� ��4��ssF��ؓI�����R T�d4�a\.@ B4��wd�:��V��òRn�a$�9$��tİ%�'�rF04��\��I�1��i(�B>���4F�o�eb@����0d��@��'2h!\g\C����� B�E��Jl�#��ˇA��k_$��0��.�:��c�ƶ��Y��Ji~�p�t(m>��r� LgP0��޵�
2i��t�j� `�v�6l�¸�ɤ�B����x��f�7�o��h�f˥41�u����:��rN0�L4FJa#]��N�*o��;#�����p�+�`Ń\82�$P�WM` SI!� @ ix���sh�$*������`�G!3��RG!�$���3�d��8�ɬ���ѳ.G&tn��b#eH\�96��357����P\UbwՋ���b��U�ʯ�/��}Ƒ#��	~U|��Lp�$4j���HVcl,)�⑄G@D2�d�(D�hAJ� �I�F# E�d��DrE���:��"�ai����e�\�K0u7������M�@���:�g��[
`U�00l74�p�$$d�ق�	g	��0��2�3���9T����	e�!��k��D��ba2���ӛ�˫pc���tbq!Ϗ���e��Q^!�	���ێ��5ä�w8M0"�]�/&2Ea�o7sI�����+b@�R�6�3�5�H0HR�����.d��U��!�����G��|���B�։@��\b�#L��8+
80@�p���c@7��t��0R,��<�0E)��`�e�qL!"�k� �!"��r�4�7��ÓR;���K�q������40$n.`H!
�t��E�Pӭ�A���ȆdL�Hi)"�0�����$H�� �lVAbb$)����:�)������(D�5�:Ƭ`
�k�8��s8�&X�A ���F�0�E\|��% A�$nMb��vx	�,�E�8�~z�c��޻�.&u������Lhv�9e�:֍��h�E��Sɯ�)]����2�2���	�� @"'�J ĆW�.�LΐѠ�	L� B�.p�m���8������r��P�М�a$r�8 +�2k&Cd>���	�F�D$j��k!5U�f �	Ͽ'8.�����}�935]��WWc���1I¸U�H�1�.9��T�`��_^�b��ʿ}����+Σ*V7��Lrbpڙ@��"���T�U�a3�L��`�2d.���`1(HCBi� U��bQ�W/� ,Z�.`����1�B�)%1��o`K�P76BKf񈆤d`�ٔ�`�I)�v2A��;M��u��#����%0����\d����!@�U4���.��)�%	t�gL��`��b��1�0eFuT�DZ������cp�#�8�0�4�8B���F�|a�:H��3��6��  p ���     m    m      	 m�       l �  �  H �             [�����     @  $   l ��m�   � �  i6�p[@A���e�  ����hi�.E�QN�k��f�@�- O۾>  mm�   �l�J�]/ZB��g��Ӳ�y`'�Zݩ�v�T @�-�,0�p�I+m��-����Kq����[VȻ`I&���٥P ����j����K2O'F�>~ž1]�J����'h�2r�;�$pkX-�����|'J�^9lN֪j8��[Y��-�����<�DK]u��J��6ث�<k<���*��9U�����N�,���aŵ6�PlS��: lT��!�q��PʵH�b�8�.:[+Z�M�U�PS��	-TQl����0c�H飭����W&�*�U��q��������*�P[VP��-�k�#i6Ӛ-[%s�mD� m�%ҫg�yQ*����B��U�y$�H����UuUJ��.��Iэ�,C�e�/;[UU$��Xm-F �K�0}���^�ߤ  [�������q�� �k�  Hph� �!mH �����bK���8ֻ9���R���9,���9R]�-�h�l H���ٰ�j��;m� ��B����>��Cv8����y[j���᪀��nj��]X�u�����   Er�  �����J��*�a����Ma.p�w[@"B�
��+�mH�j������w $�m���-m��@ke�9�ڐm�����o-@�v� m�- ��ul mHd�UU�VQڪU ��]�0^�P8�X�]�m '��UI�[��p m�����%�����^�笗�[\6��}�ײL �,�xE��-���m�
�[��*yZ��*[<-F����r���*6�l��@9�l����Xcu���������ƅ��
Z���m� -����.�M��qk���qe���f8��S:�.�fGU.��[���,�� �<��vM�n�h�[$kn��
�ڕv���Q9������Ā � �e�ۺ���۲�i �/5ֺDtU��e�9#[����@[@� H�� l��I�m��qru 6�$�SI��-� m�����7v� $  8 ô�n� ��\A��mm� pt��lm���8 ��% ���`�[@�h   Zƻq$�H}����� H ���a��.�Lԇ-� ���]�6�m�/Z �$m<t�h�   � 6��:9$�4P H �-�  6�    p   -�   -���  m�m�  ֱ�lm[� 9m   �   ���v�J h Z,�   �mH � ^�P  ���l�I� �G^��8�m� q��im  h �Ŵ6ٶ�n� p�`p   �;l��i(8�e��ۇl �  m8   6��T�SeZ�P��P   8    %��5�H6�$�mm�L���l�UU@�h��R�� �í�&��f���0[@��A�j��Iz�L�/5�G@U�[���ۖ�1�ke�m�nQ�U��]���!��Tŭݙ�,�!�p�J�*�A�U�MC��N��b�]���c�V	��3�
�U    H8۝jCk�I�ln�B@ -�m��� �  �kbm��n�]�����m7K���  ]�hݵ��@Z�)�� [N�� l�86�[���   �v��e�s�f�mֵ�rm�,���`�m [@  m6ݔ������ -�J���` ����fص�Hm��`�J�k���e[[ -��`6ر!�H��$[v���o��$i4�� �h�j��`մ &�6Ͱ�M���&�Jm[�� N��  H�SH�f���ʤ���t�ep	7k�� p�[M��Ͷ���vHm��n�6��A!��@k���Yv8I���v�V�ڳl  ͽp��zA���t��a۰H3ʤ�!��0p6��ɲ��9j�r,J���jW  �l�ۄݮ 墛 ����llz)֎'Am5��c�K$�P�R�T���+���c��E��{m��nl H$�Җ��꘰��}���r:��.�vÅ��l][UuHM-��UA �� �y�T��ҫex��)	�4:ąϪU�:%o$涣T�WWZI:lm�M� �v�Z���AZ��3���uu�����$aG�PpUE� nl�q	�&�q�P���v��{gvn���e�jۇ ��l 4��ߦ�-�m���C�I"@5V�G.�6���m������ <t��ݗX���$�UZ������j!�����-��8A6�:�l��6ݛ���P�H$��P�M�M�	��l5YYMU�cZ�۶�t�I�8 ,��l ��  	@
���T�A�+@K�;m�6ݙ m�j��%;:ݶ ���� 8H�@�L����  $ ���    ��h-��}��|	�5� ��v�  �J����$�ְ  9ml�[r��]T4��QY�@9���Ĝ| ֊ɵ��	1m #]����i ��6�  ݪM���`    մ��t�a�j��v �n�  	6Ѯ�m�	i�z�?��E� ml�t�#  m�� ��ppn���7m�l�md�����U�^Z���*�#�k��۵l�o���& � �m&o���EH�-� %�#]���8,ss�]�� ��Lv*��ضyVH�v��V���<�T��lcX'�FҊ\�|�|�i�]��=̼�W�4��<�ר�Cln4knl�k��n��		���I�i��Y
[l  �p �+�����\��7��   �-�  $����6� l �mgj$�i$�[u �	E�mհ	$NkQA��}���[l�=: ��Z   �n          �l ��M�9�� H  :@ ,�r�� 6�m�� H
嶂���6ۃm� �  8    ���6�� �� sm�6�Ͱ�vU�N<�0    D��[M�a���xh��Ku� ��KM� $8��m��'e�v��n� �m���&��i"r��'R� �$ ���`�}��    ��� J�Ԏ�~�O�m�L�!���v�i��  �ݰ������f�
U�m�	2mfs"��۪�f�vٶ�f&��.M�H mz��9��r@�[&ؐ�Z�      �9�� H��ӭ6 %�m�][V��UJEʼ�����U �v�UQNEi[���� ���6�XX�-�� �ck5@��Δ-���-��a6�   Nm��d���݀ 6��)!�kՂĄ$[p6�%�m '@v�ڢ��i�#v��Ij�[N�UmK�l�f���jkK�9٪�nڥ�*�V3���+9V`�kvN&��5a��E�4�4���dY�p
�l8�����n@j��av��Y�+UJ�m���R��L�  �`��� -��	�6�  p ����` 9#�E@���>A�  �� ݷ�@ 	J� 6�n	$   ���`m�   Im�` 	$ڶ$t]��� m� $�6ٶ��� 6�l6ͰF�h����[�r@�lz� H��Lͱ�`v��   ��  ��pn�   fu������Z� �[��$    ��E$�V�m��I��m�� l-��  x  ����rT�U��^y�Q�¼��M���U6P��[l m�@  ���@  ��hn�m6�I�ph�@ ��R`����Iu�KU6U�x<U��U_��k��{rv5*� Np�'f��"v�*�ݴJ;m��v� [P�h  ڶ  �h  ��[@�� �  6�          [x��ض�h �H���{��{��y2"�@P�1��c�O��J�~Aڢ.�t�Q�\��Pm�`DO��(m�<EH*�AGB�QX�i h�[�D��T�="0fz=K�Ph��:U���"��
�6�N���]tV&�8�P9j g���Sj�zhR��>UL�m��@�!���
�L�E:�PِS�	�pM�J8`�-J�j��Q�� l�"j+���ا
r�qX0��+`	�H�����9�P>�� �Ȣ�~~@�08(!���*c�$t ��S�	�;A6"�B��!�:Q6�pt���*�<P@:!���Qb;:S����U��=6"&C΢�� (E>q�> �~0:N�ꠅ�`!�6��h �
�#�"#ү�2
��B"0F��?<8�!�3HU1S���Q_��\��vK��ET� ��t��H�$H��m��9��0 EWB?�)� 1@b D"2�b�E"�V_5L^kƱ�g9�r��[d ��6�  p:K\݃m��-��ȢB@*dH�=lѬ�-�TU=�]�b�V��;����v��z��9�x
��ĩ���R��$��q[r�m[a4�MS�i��k�T��JY��$�-C�^��3�-ӳ���nQ4D�걛��sdu�#Ln�m]�fK�5r�Ұ�n��pY�]�>6:CEt��4�9S��Z-�d-�o_���Yo$컧���<ϡ�P��j�%D��Vd ��p��R쵔{]�aym��J�M&�u��mA�2�M�$L��`���uM����^]��R�en�l����oZ�� ʯ5A�㱜�Uj�CA찀�l�-�H���R���9�a�t�b�q��*�,����2c��R�lpQg��YSZUU]
���[��{a�N�c�ӮB�ֶq�MO&2�Iq�Ju��٪�؉}�Okl�������D @�-P�HE�[�UW(Fc"����N�GmRg�!!��f2�]�Ͳ��ml�e�v8�Ӄ8�&�ʶ�^�9y�ۭ^���և6˵�C���O�nn"��Ԕ����<���l :+%h�xN���v����ak&Yvm�j��evBT�H)w&�[N�p��P-d�[N���bc��/a�5sO-����z��5�ݶ�	
�tu�R,4��6��k��t�rێ�� ,�F��L�V����vFv�3e<�]�[T��*ҽgd��!W]M��L�*����&�U��a�R84;��]2+�@��U�T,�;Mv���v�M�JL��"�U(�8vy1nG��n�t�R�+$5J�`r�*CĈ�r:*�r��T�z�z�:��ɛn��U�mmKĻ]�d&��M؛-�jc`@����U�h[D�u�3�ʵUtQ�K 5U�H]��V��`��s���-�f�gA�75 +v�K�IN^XՁ�&�)N�i S3&s�Q�N��"(�V�$nQڠ�H!�PxlG���@z�6o89v�0w�p�����Y��M�4�huM;>y���k��ý����s���v4LvCd̦���)UAI�Hm�Î�I3�:9kU�R�ힶ�U8�*H��W=m�t\j��l3�!��a�n��b���ʬn6�*�Tٖ�u����+1�5�t���q�h4p�sX�n���מݼ8���8��6�r蹛�G��Ec��4=�4�GN&���\ZLS������6���7�<y;��O+��$"���$��P��ۀ}��T߿w������6���ԍ�NPQ5U`}�;W��؈P��wnՁ��b��v��l�Si�D�i�%�	%x���� �ژz����G��+
9+p�Z������u0>�+��3�m���^gf𳷅����}mL�n�`I+��q`=��[�KcE��UB�Yn�.ݸ"��u�Nu�!�ѓmc�l�ş'p.Y�Nԓ�(�d�J�o���?.�y��IS��Q�U�o��"��v�#&" ��y�R�����׌�/�RB\�R�R���`Ҧ~��Oߵ����0?w�7��ڣv� ��ۀ}�w^0/�x��W�	H�����n�Z���I���׌	��^x��W���p.'���#rګ����&페hMϧ�Pzػ�/7��<�4Γ][=1+����M9k��?{}� �{����� ���ŀ~���*��Y[��ՀI+�=*`}�u��+��^g&�Q��dr� ����>���a0Ȕ(�F�TH��b'�Q��8A�?}�}�������kOmM�YS��[�}��x����$�����_극�HĐ��c�+���`���ۯ主Լ����:�bҘK�n<���8��]���t>�vjqZrbn�a�JIUV��_��ŀ�ݸ߷^,����?vv96Y��Q����OJ�z�x����$����K �]n[�}�u��>��,}�w w�v��=�T�9]�8�y-X����$�������w�j�P��a�8L�&�/;�\X��YP�%r��%�������:�>�sj���`lD(Q������]�\Ak�f^��vװ=:՝�Z��ctvnlY8��^o�w����㛑6�c#.�k�U��[�V��B��A������O֦�,��G-�>���`ok���`Ҧ��{Q�D�I�V0>��`I+�=*`}�u� _ut�	)%UZ��`7��~X=*`}�u��+��d��˻8�L���`�u`jQ�ݟ��w^ڲNs�ѩ&�:��(�����)
�H 1�B���`�"E0RAp`�	� �>TG
Mٮ���5oT���b�p7�����P�\�kl�b���V�N67��ZǍn�v��hv���sE�	�uɬ-�Ҹ)]�uXgrnU�T�5gWJ<���K$���!�k�����)}�Г�s�v:3�R1���*��9�v���6���d�ڸ���R��۔��aj���%[�DkB�u`��xzڀ�8ii]�1Y�5���Yc'�*����v�rm����9z�ִ�x��ð��7Y[��(X���@#��8ܷ�n�,����;��, ����?l{���8�m��;W�dm� x���2Ձ��ݕ
�Y,���Z���� '�L����W������Y��T29V��R�{��}����������?3y�=�6�eN�9n��x����$�����,��@�n9�Sѻ��헭7f��#v��^��ub�Md��=s�s	f5n��|�_�J�OJ�}�����{V�r*9i%�j�Հw��X%�s�TI�H��&�& Œ�=p��1`ow6�݉�k��¹x�ũc ��0>��Y^0$��t�&�X�#��\�[����o������I^0	�S׶�\��9Kq�v��ow�)���� o�����\u�nGGe���E*_^��q����������ɝ��L�ب��C7n\r�\�pr䱁6K�zT�>�� �{����0��T���Sv�0;��RQ2ץX׶�����o5����,��G-���n��qjQO ���=<���u��R��\�骎l�8�[#�[�}��`M���'�L�2������jH�X�vv��	������}f[�}��Xݔ��Y-�`�V�9��Tn��F�x�f�"�U2����K[N���Œ<�F"�`�vY�wn }�[p��� ��ݘ��m�"��]j�*����(Jd`9Ǽ��:�&��?E�$NWc�'�j� ���,o��=*`Y�0/����q�e���V�ȗ&�� o����h�»�!(��:�ڰ1��|Dqf�%��\��OJ�ޥL���� ��l��Z�:B���[�ﹾ�Q��k���>K���ܹ���\�/nm���g^N*��-V�G-��|z�ow���0��� ��U�Zq��[��&�����@��R)�����}� ���~�w >�;�j��ܪ�3�,`M�� ��0�n��W�݋�=�FQ�Ѵ� ;��p�n�X��ŀ��}���t�6����F-��I���׌��d��;��p�ȅ�)����Q�Z�-�(��3�\�*�F�]�F�yK�ݢ��%7�ǭ�v�Qځ�$����Iu��KApa�uHϹ�&&�<tc����2�s�M���?մUGC�G�!#j��z��,�h��2X��]�u��R��7l$��}��q�u�w3��p��Z_ݨr蔟Xlf�P�	Gs�!&ݺx�&�'L�*:/�Ms��] �����w�>E���\M<�u�=mɰ��Pu۫O�^-����M���e^�H��1�!�]]��ذ��f w�v�~�x����,r��	e���%�=*`}�u��+��X�#��-��e���ۀ}�u����M����w� ����P얩o���K�[^0=�^`J��m�+N8�v��Xۻ� �fN��|m��z]x���^kx��\]��ضb2��lf&^��p-��xw:R����VαP7\���l{d��=%L������������=�����-N�0�{�* �BP@����3��Vzݫ��� զ�l�2�WZ�[�w�tŀ}-x���y�I*`z��˝ݛ��MӰ7�������e�$��=�1`n�e`�W KmX��X�Ky����KVmڰ5(����{����Uv&�f�������G�rzX�kok��:H0;:�jLXU���λ<�v2\��?o�߹�=(�m��/0>f��m��%�[+����V,�9�&�{�ŀu�}0{�0˦�9����mC��ww��va���{��e3����H�1��֪.�CqP��]1.�:ܲ � 1���A!$H�
�8D��Ca���A�d`F!��3Ph�#$`�Ϧpxg�N�iN���w�5ے�R�4�Û�2�
!U�v�Ev���U�
"��r#��
�^�Í3D*�|�z�Pv��"��S�E0���s��vO��M�����ܪ�E,��>�o� nﯸ��x��a�9�{�`k�kjiqQ'*���˘����,���~��0=�Y�$���g�F�md���p���g"ȗ�N�����,rpl�lv�c�����mR��nWZ�G-�o��X��o�_����͛�������/)"nX���)X׶��K���o�ϔ)�^��w�X��>a�޾r�jK%���V�(S��́�Q	Kǵ���Ձ�ǋ �����D����ex��ۀ>��X<v�%u, !@�	(�P�ƬlACh�_�����]I>���"vT��jr[�o�� ��f��׀u�����~��啡:쉢oT��zFNٰ���3�Vi��\s��G�8�խ��]���q�붢¬ �{� ���`]���Q����q��[��wiܓΗXl����x�-�07�7յ�-\����0��<`ʘt���뻊�Y١��U��W,�e� oY�:��l�{<�aݏ�yI婰����M�wj��ǳ�G�;��}'b|������K��#��֫��K^9j�׷�/4�駥3L���&gs1�ۨl
C�;����">`n�q���d�iB=��=T�n�析�a�<�0���3�;L�Q�)���E���s��c�v�Kvi�8�T�!�;�6���N�z�S����0��o/4ҹ�ݔ� ����o�����ې�.l�W4�;���;v;r5���ܮc4��z��]k��1�{����/#U���5��m�m��mM�sۣ��	���˦���Y�ݖ�r"�1��$���% �����o0/�ǌ۷ �����DP����{�0�q� �������KL���7�rY�#�����[j`Y��^����h��Q��ڋ
�v������o0/�0.O���;K�-��w^�wf��V, �ݸ��A�`���%���in�7�X��R}�n�۴>�8m��V�{4Nx.�F�-5or��o0/�ǌ[W����o��|2�:��ƭ�[0�j��%B�	BJ��{�V������ٞ�gv?E�$c����U`�ڰsٱ
e����Q��굀{޾r�i���
�n��׀M����x�%�0>��;;���%��\��6��	�G�[S۽ـ~{�ɱZ��1�Z�j�Y/;�˷m�\Z�:mK�N�v�\tq�ĥ�q"Y�nܖrH乁=(�Kj`{l����ـ~�Qͅ�u�QaV wmLm��m����x��?�\f+*v��8��ـu�����+��4�g(�Dr��s��ѩ$���u!�����8��k� ��ـw�tx�%�0=�^`O�M+B���b�r��\�3��V������:��=ݘ���č�j��r��C�T���F�F�ެ.�<����d�vz2b�y{V���*�}�\����:�v`��1`�u���,�V����x�`d��`g[V�u�(�:�ydN
��$[,�5�ޘn�Xy.$�f�޸_�� ����'eNY-R�Kf��������z���fjX	"�` ���#@G8�q{��������D�G$v�&�+ �7V�s^��2u�,�j���ޥ��5�)dHa(;��{m�(;��;;Ev�]����ݬ�$���]����L��USɪ�����X���u�ka|���� ��ޯ[V�1�f��|�y$��_��X�z����#͘���+����V, ��ۀ~{ݘ�ـ~��-Q�R��)�n,`֦���m������n�X5%���B�ۀ~{ݘ�]�{πy��Xu��dQ	��r]��4E�^�������a�s����m���m=�H��i�X�,9��j(F��hc9yV���;i�BNJ�nC������Y�8�6	�`nLmkh�x�J����'d$���	��m���ɮ��s�q�k��j�g!�m�gT��[�==�i�t�E��m;��.8��^c/TWg���m��������du�S*o��s�#BU�-�����{����v���(W&̽;�kc�n��cqֻS��FZ1�o�<��n��[<;�˳��|��r�ζ�Xu���N������'eNY-R�If�۫!���IH���#����o_��cm��{��o�6	�A�$��ڇU�6�}��~���my�ww}�^�������������eυe��;o�6�^�)���M�Ͼm��Ր��o��o�6��M��눭K��Y�ww}�^����������Һ}����qLm����3m�����!�k�����5�2\u�}���v�C�]\.�u����,e�QX�`��Y�ͷٺ��o��4������1�����ͷ�cرE"-�dą�L�j�o>�{w���6�`��r^*�o���ƭ��s����{�| ~?~���`{QG�����1�������.I6{�!�����|����&�crR@��K���~���ogud1���ۚ}�oˉr?nx��o��~"��,��lnW�ͷ����o������~������u��m����?}i���my�n�lg��u�m��ɼ�]v1�����K!w����U�U�u�ۻ�$t���ݱU�ww}�n���v���߆�6���s���Gm$-��6��ݳ~��Qʪ�[�z~�fg���s33޻g�zH����늎Yav׍��;�c{����hƭ� hth!������m�o���}�tfϕQX�`��Y�Ϳ����~Sm��x���{۵�oܓ������ݯ�b������*��o���>���=���m��w޿|�z�LSm����~$���hZDՊ:���DӧiRz�d��/i%z,OD�mI����ú�Y����~��o�}^6�~ݿ|�z�LS�H��w<}�m������IGZ�Z�ww~���fwvݴy�wwd��}��~�/�� ��o��=��r�M8��n�<绻��t���ݱU�www�Z��u��Or�$v�XU1�����>��oy���[m���w�n���ad�  E��I		�����$�V0&��z_�Cm����Nڂ�-��6�m�9���?�����ݝ(�{��=]?? ?������z��p4�u�2<�J]�Wq���u��M4%Y2s�:�n�9e��Lm��ov��m�wL�6����y$�~��~�)�������ʪ�b�RI-������I%�ks��|�z��Sm��v��m���,QH��㔰��{�sO�m���S�9�r����6���cm����
���Y[�v�}�m�n�1����߾m���co�I���|�}~��&�c�+"l�ǻ��J��wvl��{��lt���ݱU��n_��@2)Fφ+ ��BS��a�D��#��i
��p�!2!�ؒH,0JGY��A�	��$�03�$$dHĐ$���,T�# ��0r�=����/�"F0���b�#�YQ�� �cHF1 �Xb�FB�3�OA��� �C�Q4h��$0eM �Ñc!��cQ���4	l��J���ЁD��� "��P�BH�b�dd$$FH�N���`�A!F1a��FA�X%d!���I3���p�4�bJ⌃!��1dbB)ÇG�{���� Ĕ�n�C��*:�n�#��e0!i�DL�	D�, Cn���b��D C<,	$T!�0�X� �)$H�$�H�"1 Abk�8%Ȇq��_R����b0	�@"4���:��l�m��$մ�gl Z����-���H-��L5�ZD�[�-�	��v8�툪q4dv�ۭq���t��s\dv�
���\ZB9�\gn]֋����Ʋ�v��Yg\4)*�ӦQ�w,dM�/���l8y`iƉ�jۮٲ���/�rP7lv��K��ljn4����-D�#WmT�X;Pl��T#c�*�,E�܋.���*@�����-��8�$�/J��k��ZLu<��m�<����6+���pX�G�6��؇�������Vaղ�FÎuS��L �UR�2g�r/r�Ή`���^Q�Z�D�Լ�r��j�ns����IC���9�erҭ�ӭ����(kb�k6�U]y��6��iz]6-�������γ�x#S��p��v��G"�<@�J1����G/;�mX��Wm���\l5*����H���p�N��6E������m�J���UjU��WC���a3��Q\ŁQ�2m���;hyܩ��g)l�]�_F#t��7@�ßI��k�''GvL��[T�ݠ�.���tez�v��SܱG`{n�62#Q��ض���ɪ6/' � FʍPSU�8Ԫ����t%���iwI�̝;"O[uAȍ6�jj�7l�sPc�pN��*`�<�5�mg����H%I�˶��W=`�W�WL���+��-��h�ki��Si<�Me����c����˵*һs��[T�&n��Z��eZ�gieM��@
�ڰ8���᧊D�d�c�j���`V{gk� ��+�Ҕ�
�B���~U�hN�����������v�9eYqp򩣬)��۲���y�y�N^��e��0�,g��f|��Z��nMJ�[T�UA���,�`��e`��U�vB�u�?|l�̫U.챍W)2���ULuplѻJ��ܩ��-���X��l˥��fz&�%�:L��U�\���` sv�\��*&�u��M �|��(�b*tplt�!���N���!!:�Avl��kM4�OMΆ��z�q�h�F���'I�^��	�v����vsŬ��v ����b�	=����3��i3Z�몲k���.��6��pk�R�:+��둔�4�i�F�y�m������`d��]C6��b�*1��<mft�p ������?)�=I�����l��k��ڗ�6��s˘L��[�:}���84���3v���q�|�����$��K�p��۞[]E˂��ڠ�k��nIjg�������<绻��O��ݝk�����/}��￶��A�$��؋
�6���i���\RG���cm���_�m���cm���wC�G$�֜��}�m�n�1����o�?s�RM{���{��K�����o�-��G-���a����}~�����)�����>���7r�o�7G�|���+#�߾m���cm��sO�m���^0�����? ?D�"�G�[����tk��!^��;���t�ŷWfb5ū���z祩��r�Lm���i�Ͷ��k��o�ݿ|�z�LSm����j;%���8����u��iU�a�(D��dCL&a�(�j$�u�W�n�ݔy�wwe��}��3;�f�����IIe�6�{�������<绻��O��ݝk�����&Ӿ�eU�-��ܷ�o��b��o����o�w!��.%$�o��6�y�'셎9�Lm���i�ͷٻ���o�ݿ|�}}��������+d#�2�bً<�3+Ӻ�Ë!�;x��[/1�sGE��''3NZ�e�������d1����_}33����BI/%ک��m��陟z��{�A�H�g| ��������e���.ff^���fs�����eǼO�|���+#�߾m�?�6���4�w�B0%u��q﵉�m��ﳽ�oq݋��j((����o����������o�{�!���w�~�������V������Ij3ئߟ��� ~��w�~m��=��m��sO�m�Ӈl�{�j�*�H�<��[vL�[<��r�mrp�A��rud��+������ǙE��u2|�m���l����o������ѷ��cm���'-U�-��ܷ�l���䤍�<}�m�o��m�{��$}稽���!c��e��{��|�{;�o�G��_�m�����m���wC�"Z6����~�����}w�m�w7�:��&��j�	B!sA���w��o��ޘ�q��#������o�ݿ|�g�]��}��|�{;�m��ZƁ�ld��)3B3�
�uz�4@$�mqة��u�a��7]t���-~~ o��?K��:}���ey�wwvYW�n�ݗ��rڥ��NZ��o���Ｄ��}�c}���z��n�pU4K���C�^0	eL�v��Q���f�5K��"ʰ�ݸ�멁,T`[+����.�䒮L�*���Ձ��ޟ��ՀcǝI*a'�y(�
L�d�>=frru�frj��nȹ{w8�=c[��K���p�	�a�v�u�gs�����L:�;��Ǭ�δ�l�X�2���c[X�$Apő�ۮ

���������-� �j�="�=ѩħ^v�h{d��+��rv6���f����}o��T���خZpn�p系��"����v�h�k)�ς8,NIqR�0���9�&�����-�K¸�D��֭ێG8.�`wi�Uέq�g���;oj��;�o�".�F���̭,�ڰx�����ڰ:�k�0E�;Hղ�`��Y�&�}���|�p�n���ީ�G�v�0	eL�v��Q�,�`�餘���t�X� >�Q�,�����<��R�1vorԘ�F��`ʘ�^� ��M�E���#���ȝA�n�ܶ���y=5�L���\*�n"���n'"+C��I䅝���`_EF,��zͩ���� ��viP��(�%�� ;��u�6EY�@�,��Τ����o��3ˉqq�۠�[T��m���LO��0'��z*0YS�?h��,q�+-d�ۀw��0�ۦ ~����}�Pk�0E�;NJ���,�S,Js^���v���0��=�YA�r�]��:�{f��6M�-��V
7`�v��8��M��W<�G�����Z��=eL�mL	b�v�~[��bj�Gb�H� ?nK�؈J!)��,�ZX<u`|�b��j��U@rWn��� �ݺ3��س;<��|��mL�WxA�ڵ!,Xr\��T`ʘ�ڰ=��'���u�g����G-uYS ��SX������������|��\4t]��7W;�˷m�F�^t�n�d���:8�d�.Gm�J→]������Ɂ,T`_EF,� ���'�r
�Y-v���0��%�0Y�0>�nk�g.[ۉrH`_EF,��zͩ�7�L��oa����eX\�92��X^�Ձ�)�
)(��Zˈ�9�����zi2�[,U����ژ�F�T`ʘ������6:Ҝa�ZGmz�a9�G�C�s���ld{b����B�9��v띅�/����0/�� �T�=f�����SQ�ij���`��L ��ۀ�kۀw��0��͌|�G%D����:�Հw�]Y�D(�2�kK{���������ۖ��۵0'��z*0YS�ަm|.���%�%�0'���*0YS ��{p$��qw�["�	 ���.k���I�Ƹ�����D�6�璹-�r�׹	������CT�m�Y*��p;[VtN��e;t��v�g���2\�C���VU�Iy؇�۶��[�p�I�Ͳ\mi�8��v[l1xۭ���9؍ƃ���NbM�
l�zƳq��9�kh��'V�of�q�����.��v5��6v��"te�d�y.� �e�]��W店��G��Zꔲ$*��b����9w����=/��m�i�D`k[<<ݴ<Z�W��I#�?H��=eL�m�m� ����eq�G-��]� zʘ�ژ�Q�})v�(�*ԎKp����;�n���� ?ov�n�X���Z�T%i0'���*0YS�f��w�`~���MGl��Q%��7�n��z��;�.��X	,f�#~&�r�[�����Ӻ�v<q�BuX��v����ju�zx���<I����o��$VD;]������z�L	�����`��-XA�m��n ~��n%�qq.�~��>�F�Q�K*`{��ͯ����b��Z��׌	����ۤ��&'���>��XF�N��Um� ���0�n��r��aD�{�;��v�UI9\��v��wn�%�z|w}� �ݺ`�{Fm��o��i�e+�:������)w��9[�녮�<�en��������Kc���#�߀��=0����1��""�� �������+S�U.Ua�8�.`zJ�}�����6g���޾pU8;ev�	-X���jI7��:�ع������y�jS*Dp[~���)��d.7D5��|!�)�&8���WC � ���a#�fwJ���&�55�D�xd1d�����)�G;W+~���� �&&0(d�ϝ}�M�u\�QAڪ}C�%o��T�B��U*!�x�G �E٠ �����'����b�??�&��Y$�Ȇ[*��}��&����Y^0%���P7i�E��ۖ��ـ{��|�}�ŀ��p��$��8[�ny�r���qLx4iƶ���=\s�l�؞7/W]�d�*d��`u^NX:�VZ봳�;��,�W�z���췘L	��۫�W��o%�Y^0	�So��`zˋ ����+U���,pvU���p���f��k�Vk�VWL|���U��v-���I�/L�����Y^0���n�wv,N
�-B������W�	ex���y�/L������w7����1q;j����Oq�ty��M�Ǭ���"ܫȝst�xi�u�%QN�Mw�����<`M�����X��`{}��%�H��d������?wn� ���X����>��7�LUr�hܳ ��������׌	�XXf�A�䂶�I*0<���� ��ذ	�X�\L	��ڻ�\,�guR�;�ڰ6Y��?�kQ`w�ڹ&�3Z�� )#TLaQ�AU�@`Ȑ)�$E�B��� P �T��M%� �\�����rJZ�ӎ�kH��a��ɻx�ѹIy�1�F*9\h.��d���:ܶ���7'g�����ư���]��uX�w&�T�뮶������g���M5�n��#��Ӳv֛Gn3���.��6%0n���m��M��Ӣ���FĆ�v�Jȯ�pim�����s�8w4�3eًl��ǰ�i��<Ԏ��C��xܪ�7iYynl�ū�qD�h����֊Eb!�f���L��W���v�P�`k��]�\�g:�뫭M�Z���Yc����=� �ݺ��k���<K�H�x]�s��Z������n�V��k���^�݋����^DT`�n��;�ڳС/˜��zl�5zl�ӞGm�� � ��q`~�� �έxO��|��x�M�Y$�ȆK*�>��S�kg�3ڰ1�`�Y�kT��U�%���d���ڭ��|�n�{s�mr�v�ۛj�N�n�j�ʟ�z�ٰ;�v�x�yG��n��=�~�:ܐV�Ӑ� ����*p�-~Y�
KЗz{;�V�=�`c�5���5�v@v�'mXw�� ��nl�
e�f���Հ�)�u*�9\��%X��w<P7�O<�ݪ��'����.�酤��X�Q�.�'�����`}ex��u����~�O��M<p��P�j��^yK�{t���㭺����L��K=���v��w�|���ޕ������C�K�����V���Kk�V���,���=*`zJ����?m�囿�wl���Հ~{�L�?wn��b�J 2D �(ED,D�V(h��Pv������ԓ��jI�9 �H�T1�m��f���� ��`~�Ł�>�o��{D���I!Ik�.I�=U��?~�>o�����Ϳ��v����[hp\��%,�NJ�0�7N�.��v6����y'[f�VWkZ%ؠ�Ԓ��`{d��>�������� ��o�Z���Yc�r���vg��z�������+���ŋ��@���ԓ �Z��Q��e��0�p��'j��^D۶�./����ŀ�}j�3�Շ�[SU.�X��,��U,�)�~�w��޿ ~�z���L6�(��-N�s.���u�=��U�k��m�8��l�srig2y\ˎ���������޸��0=b�ޕ�����7�In�I�}�S���O������=�s��l�{D���I!I+q�p�|��J�OZ��T��;�zW�
;eX�O{��`��� >�����}��wɿaJ���8U`}8�,(����n��3��X��_�"�}$Q}��G�H�E[1�NZҺ��ۘ۲�p۶n״��4��ÜmGn�:m�wWH8���]�p�<��
s�vҦ�+� ]�݂�H�ۮM�!1�,,�oC^ydql��һ�Aq�F�Ƹ9R�z���%9�t!�>tq��8�r�e�8��K�H��n�Z�cX�a,C�����p�6���]������;��s�^l\/n����������`��'aݦL��O�յ����cW�qmr��qg��k�jK�!�;�,����n�ֹ)��K�����Ҽ`}��`_K��JKP�"n�p���?�.qq)�Ł���,��W�%&g�\	���{�rIO����e��=�S�{t�>�������Ki��s����w���X̦Xz�%���Ł���I1J���$�`��n��T`}*���l�g^�o%���&pPG/Z�lp��]pK��X�t�J�t�'E��h�<�8�$�������;�ZXc�Xu��H�Ձ�����W�
;m0��L�.u%��pI(�J-��VS� �qՁה�ԡK7|����+�:�� 7���ݕ0=ex��UF޷��$j�aD�UV�S8�Ձ��Ձ�:e���7������X�-rȚ���m�?n;V�.��> y�V��V��R��]Xz���v�KۗF��α�f��n6)��7���NT�{���_t�Y��[e$��=/� ��0IS�W��{���uKi���s��a�{Vk�V�闩Dɚ���9k��G-��-���\���Z��\��D(�DB�s����[��pR�ӒB�V�-��}���~��� ��ہ��\�{��{ux�S���	������e��^n�����)�������@�7`���V��\n���6�3�k��p@�-�p͒�%��w����@���ڷ�$��,��0	%LX����� ���
���yb�Xݷ ;���B^����kŁ��x��u`}����euX�S� ���`n�0�l��� 7w� ���`:J�R������ޖ �v�3XW�"i�bV �8p6� �/u�@k��Q5K$���)m0��n�	z9�������`>�e��ɉ�U)�+W8�ZC����9}{I�^:Z��n���nx��}6r�vnn$j���o������v��Lߤ��`8�)��52E+��In�{���.Ho��0���p{ݹ��8�=��HC���v�J�����3�՞Q2k{Vk�V�Sz���r�d��`.%���޶��Xx�XyN�ޖsw����Wn/�ط4I&d���+��Ta'>�s�$����,H�5r�r):�@����DG�|��C*�X� �ω�9�K�4!G�T¼ "	4�Z�㐴f�,l�P>�D�G1�&B4"1Z��Ta��""�p#��s�<��E�H$aT*�O���@q@�  ���\E��EBm�c�ٰ8<D�����+#��aA �p������������hG�!�\�L&�3�(F)����9ė�$$A$��9[�"��m��	 ��Jj�m�� Zv���������+j�\��Xň����6�[Kj�WYY�^�՜�Ǔ��$�
��n�n7Xv��dyFR��l-����ӹ�h���/2�z�M8ȸփ�]�y^�\�!2����R�흀�^낋���z`w[U�f�xव�-i�$�ְD�r4�y�P�Z�k�L^��Xmr�&�qȏs���j��v+�u��ێѬ��P�]�磷A���b���3�}�X�㵻 la�mɻvU�n[n�j˱�����5UO+�R��9���a#e�Ć�g26�u����6���ӡ�#KTڥeW���q���UU*�N��P*��@<�ם56�.����G��H[��[@�Kf�,�k|D�OZ�t6�nq��.y�7c�[�#'�E�,'6;0S+�"1{crG6;pm:��ؕpH+j󶩻U)�F2�BE��LD���u�j�p�B�:W6�j˄��m�I鉩�-T�d�����f���<�N��\��b�g9��u�`�s�9G)�v6�gk҃�� �u1\0gh��&� H[2��V��v:��4�5ө�M�tm�q��S�r �ԡX�ڨ)��yYY�j��������e3β9׍;D����F\jj�Ǳr�t�ŴJ�n�6�ur�AJPj�K�U��F��Y�kp����V�[Q�RHxVGIr�!=M����췝�;F���F�UJ�R�+��N�e"ZU��D�ʵr��961Ҫ���u���o�ҺK;P�жJ@9jnn���l��񐄭�8rH��:���U���Fegv���3�������*ԥ��r��i��쁩q�+��̱�g��z�ׅ�ͫ�GC�%�"j�<����UpW-V�ڕj�V�R�@5*�TpY�UiV��ڕ�Ŵ/PXֆ�6Z�i2�:�y�'mm2*�FY�Ӹ٦b���Uff��N�g��c��f ݵ�����{�������G*�T\j��P2�h� �A؏���p��d�"�����Yɓ���gٮJL�����(�����s1٭�;cZf�9��9��Y��}���S=p����4��W.��W;�w�͓�'tmp6rfk���W�bӵ)ĂnN87xѺzv���G-��u>��&�#�{\�]�\�)��p�`�v�A�(q�S���9�3�;rC.�s�>�Gn9�m詵9��mm�0c�y�&t챐/����Pj����a�:Du1�q�����G�ð��ϋA�4�my���Ź<�)U����;�mX��`���0=��~f�?!�VXV@vʰ�T`֦d���+��eYٿܻ�yoq�$�=j`������L���1J��[m��n��{Vk�Vu�,6&^nՀ��إ�8�rV����� ��`z�X^:�<���C�W+W(�q"�mc:ع�u�9õ�>z�h��E�ݴ�XF8�v��*HB�e	+vʾ{�� ;�v������q`��e��*��ns��$���u��"��I������z�?��������$��EqT�*��5�Xx�Y闛ZX�޸߻�-qѲD+ʛv����������0	�S �T��Isn���(Pvʰ��L�q����{ݸ������h�9E,-B,*����s��;^;c��걎�mh.K�ٶy�x����8��<�,���$-��8��޹����&%�y��:Mı,K��h?$�&"X�'��_��q,K���I\o3�[m��nq|q3��L�}�����bX��}�I��%�bw�צ�q,Kľ罝&�ؖ%�ם���3�����l��s��Kı=��f�q,K��=�M&�X���1(���~�15���gI��%�b_��q|q3��L����!�����Yq�I��%�� b'����q,KĿ���t��bX�%���7ı,Ow�٤�Kı;��s9�&n3��c79��n%�bX������Kİo=�gI��%�b{���&�X�%��{^�Mı,K����q.3��J/�89�Nm��#u�0{Na�Ρ�؝��\�x�[$q��9z������=�{�K�w��n%�bX��}�I��%�bw�צ�q,Kľ罝&�X�#8�w}��F�#��*�v����g8X��}�I��%�bw�צ�q,Kľ罝&�X�%�y��:M����&qv�O�n��b��*�/�&p�,Ow��M&�X�%�}�{:Mı�1���gI��%�b~��l�|q3��L��7g����9]����-ı,K���t��bX�%���7ı,Ow�٤�K��X!#��"|��}����I��%�bw���ԕ;��[�����g8�����t��bX�'��l�n%�bX����Kı/��gI��%�b���q)����'�X�Y�9ej�	9��{t��û7d�!�p�{\l��B�� ���y|_:�8�r�G-�/�8���/�{?����bX�'y�zi7ı,K�{��n%�bX��ﳤ�Kı9óؘ�-��V��g�8���-��q|�D`&"b%�w���7ı,K����&�X�%���^�Mı,K8��M����r�d��g�8���_s�Γq,Kļ罝&�XbX��u��Kı9�k�I��%�g���[+U+Ui�ۜ_L�g�y�{:Mı,K��4��bX�'9�zi7İ�/y�gI��%8����גּEXH�B��-�/�&qX�'��zi7ı,Ns���n%�bX������Kı/9�gI��%�bAj�z� �O`�0\�.�C'�v[�x��G6w/��C�.3n'�1���V8��q�tl]����4U��]�v��.+����-vʝ��ۘwm�n��UK)���M*�t	�V��'õi�^���5� �8y�X��z�|����1D���cs��q���ֳt���)�N�MI�;m6���6����w:t�N�9=2�È�K&�9l�$r������W�������/;�����˶�gm�V���h}=�[u���;7��v�Ȝ��S�k%u�^��YۘO�ߤKı;��zMı,K���t��bX�%�=��?O�b%�b~����/�&q3��^��?��%����\gI��%�b_s�Γp� �LD�/{��t��bX�'�{_��q,K��=��7Kı9��}q��d���s��6�9Γq,Kļ罝&�X�%���^�Mı�ű9�{)�$�Os�Δ�I�8��[.!q-��j	 ��u��Kı9�{zMı,K���t��bX�%���7�L�gz���KhJV���g��bX�罽&�X�%������Kı/=�gI��%�b{�צ�qL�g8�Э�ҖZ�a]�duږ���l�f���:Mu�I3��c�۵�a#m痫���\��+���8���'���8�8��%�y��:Mı,K��4�H�D�K��~ޓq,K��[�[+U+Ui�ۜ_L�g8�}���p���dLı=���I��%�b}�{f�q,Kľ罝&�%8�����lab�
�ݷ8�8��bX��u��Kı;�{f�q,Kľ罝&�X�%�y��:Mı��/��&��Zʭ��8�8���,N��٤�Kı/��gI��%�b^{�Γq,K��{�M&�Y��&q~���9lnJ[!eY����%�}�{:Mı,K���t��bX�'=�zi7ı,N��٤�K�&q5Ӭ�ΖZ�)`[U�c�}�W;y�׎6wL7vv�9��zض���q[�Y�F锱�m��m�����&q3�����q|qX�%��w^�Mı,K���i7ı,K�{��n%�bX�{��x�ŎJԵ��s�㉜L�g}��8����q,Ow��Mı�a���}�߳��Kı/{�t���Fb&"3�ux���)m	B��m3�㉜L�b{���i7ı,K�{��n%����8����7�_~Γq,K������Kı;���s����.q���3I��%�b^��Γq,Kļ�}�&�X�%��w^�Mı,=���4��bX�';�u'���C93K3��I��%�b^{�Γq,K�绯M&�X�%��{�4��bX�%�=��7ı,Ovf^���i��i��K�]����P=�.�lvqm�Y9��C"�Q�q=���*�����%�bs�צ�q,K��=�Mı,K���t;�bX�%���7�L�g�o�^L-eV���i�_,K��=�M���D�K���gI��%�b^����7ı,N{��__˜D8���.���(�d$�ى�d�n%�bX����:Mı,K���t��bX�'=�zi7ı,M��q|q3��L��=��Wc��sn3��7ı���t��bX�'=�zi7ı,N����n%�`~��#���MȚֿo:Mı,KϽ���,q�Z��9nq|q3��L��^�Mı,K�����I�Kı/���t��bX�%���7ı,�~��o������;(�W\Y�
5ma��wI� 7g/ozD��wX��S��������6�9�Mı,K���4��bX�%�=��7ı,K�w�Щ��%�bs�צ�q,K���K|o9�Ì�����s4��bX�%�=��7ı,Nc��4��bX�'=�zi7ı,N����n'�Ab."b%����G���Z�L�����g8�ų���I��%�bs�צ�q,1=���4��bX�%�~Γq,K����i؊
!�fq|q3��$��u��Kı;�k�I��%�b^��Γq,K�	1�����n%��&qv�M&�ұD��/�&p�,N����n%�bX+{�{:Mı,K��}�&�X�%��w^�MĤ)!IДy/)��OnyER
�METu�nE�1^��P�wEn8�s��1�;>.ͽ\4���E�H�M�Ae��s�=X�K	���a�rOj��Lb2i�cv�������)�1��V�:�ϊ!�khF�7\J�	(չ�lupc�ϔ8�nn�ҩv�C��LP �lg��e5ųl�V�<����&^��`5��c��2���@b�s)6��:����Z�9�s�|#?8��e��-vZ�\�C�{��;R���s[�m�!���
�q��R��D���d-��~8���&q?��{:Mı,K��}�&�X�%��w^�wı,N����n%�bX���z�8�r�mn[s�㉜L�gq��Mı,K��4��bX�'y�zi7ı,K�{��n"�bS�V����9+R�l�����g8�N{���n%�bX����Kĳ�{��gI�Kı;����&�X�q3����'��Ptv�-3�㉉bX����Kı/y�gI��%�bsﱤ�K�V�绯M&���&q{�i�/��rR�d��g�ı/y�gI��%�bsﱤ�Kı9���I��%�bw�צ�qL�g8��q���2X��z�m���!�
�n����ƃ����Vg�ً�~�w_!�j�Ö��-�8�8���&qv{}3��X�%��w^�Mı,K���4�@�D�Kľ����n%�bX�￾V��b((������&q19���I�l
���N�>D a'��}Q,O��zi7ı,K�w��n%�bX�ǻ�i7�*b%��{�5��Zʭ�U�_L�g8{���i7ı,K�{��n%�bX�ǻ�i7ı,N{�٤�Kı_�u��+!%��[L���g8�����t��bX�'1��Mı,K��i7İlN����n%�bX��P�	���mn[s�㉜L�bsﱤ�Kİ��1��~��}ı,Ow��M&�X�%�{�{:Mĳ��L��݊zJ;h�J��[[��5�vō��\�(�(�Z�j �D�*�tE!�i�;���m��%�8�8���&qw��q}ı,N����n%�bX��=�i7ı,Nc��4��bX�'N{�X룀���Y����&q3�w��8��D�K�����n%�bX���߱��Kı9��f�q,K���F���9�J풻i�_L�g8�w�Ɠq,K��=�cI��4_�ŵL� ����
k��Y�(j�(A� ``$C)��?|�MdQ�$B3 A��& p��@Y�(&*�I �V!F+CG(T���rB#@�	F��U~%2e i����@)��b�@HE1(e4�U�]���j?�6�Kk/1�6�h(|}Q�`�������t>]� 	�2�誡TTҽQ.�:S�(���1�5�}�I��%�b{�צ�q,K��'m�=��Ŏ0f�9�4��bY�H8�����Mı,K���f�q,K��}�M&�X�%��sޙ����&q3��w�*�N��Es8�n%�bX��}�I��%�a������%�b{��Mı,Jqv{ޙ����&q3����X���f�<�n�wnmڵ�r�-nk��a�,8p��l�I
H���д/"vʳ�㉜L�;�k�I��%�bw����Kı9�{�Л�bX�'=�l�n%�b����s�O��IcVB�g�8����9�cI��%�bs����Kı9��f�q,K��}�M&�%�L��Џ�l���G-�����&%��{�Ɠq,K���Mı,K���4��bX�'q�{Mı,�g��?}v�K�K3�㉜L�9��f�q,K��}�M&�X�%��s�Ɠq,K����U��xx'3�~�t��bX����/�,�@U�v����g8�O{���n%�bX��=�i7ı,K����n%�bX��}�I��%��/�q.$����9?:�7xGm�M�PX��j��[����p���V;�|����%+�J�q~8���&qzo����Kı/��gI��%�bs���&�X�%��{^�Mı,K�캇��H�|vٜ_L�g8��޹Ÿ ؖ%��w�4��bX�'��zi7ı,N��4��bX�'��Z^*Ъc���8���.�}��n%�bX����K Fı;�{��n%�bX������Kı>��x�g6dɗ�q�I��%�b{�צ�q,K��9�cI��%�b_w�Γq,KP�9��f�q,K�]���
BK��8�8���+���t��bX��B8��߳��%�bX����4��bX�'��zi7�L�g�KW4_�|��m�����u��)3�71�p��ƶ����+ڮ�Y�0t`�l�hUۇ��ۅ�K�`����؃[uN�f���C��{vĒ�-���ѩrWf�v;p1�EX�bi�;�p�q��=in�a�D��ۥ¸��WA�v�%k�����6��WnU]�������hq��:���3��9#�7A�݀�j�=�M��',���^�d���{��q{��v~��AuG�D�y�={m�W�.�t���0����`�.�;���Mۧ/��m��s��8���'����_D�,K��i7ı,Ow���n%�bX������Kı:w���,q�E,u�-�/�&q3��]���_D�,K���4���b%�b_w���7ı,K�߿gI������$8���?��>��\]j�/�&p�,O����I��%�b^��Γq,C1�����n%�bX����4��N&q3�}�7����JWl��L���q,Ľ罝&�X�%�}�{:Mı,K��i7ı,Ow���|q3��L��tx�9"��[nq}ı,K����n%�bX�=�l�n%�bX����Kı/y�\���g8���o�č�j�j[	 ntbѷ=N�q�9��޺xx�Iv���Ht��V�(;h��-�/�&q3��]��f�q,K��}�M&�X�%�{�{:��&"X�%��߳��Kı9���?f�L�2��s4��bX�'��zi7�&��
�&"X�����n%�bX������Kħ}��8�8���&q{w#��G���.fs���Kı/y�gI��%�b_w�Γq,TK�绯M&�X�%���^�Mı,K��=�q����g�&s��I��%�b_w�Γq,K�绯M&�X�%���^�Mı,lN��4��bX�'N���&qqm��:ݖ��8���.�s�q|q1,K���4��bX�'q�{Mı,K���t��bX�'z�����/�vu�B�\���c��=b�>S��v��Ѝ�������4���o�ߛ�D�,Ow���n%�bX��=�i7ı,K���Ю�X�%��w^�M�3��L��kM�}ls���v�8�8X�%��s�Ɠq,Kľ｝&�X�%��w^�Mı,K���4�����&qw�<<�b�H4�8�ı,K����n%�bX��u��Kh��5Q=�k�I��%�bz{ޙ����&q3��w�+J���P���9�n%�b���^�Mı,K���4��bX�'��{Mı,�!s��U���$)!I8{į)*h(ɗq��i7ı,Ow���n%�bX��=�i7ı,K����n%�bX��u��Kı?
{޴����K���n"�qc^��F�=;%[۝�hV�g���"��<I���,�k��IE-���,K��1���Ɠq,Kľ｝&�X�%���^�Mı,K���3�㉜L�gwS~	>v�2�evۤ�Kı/��gI�%�bX��u��Kı=�k�I��%�b_s޹����J>(q3������8�:�q��7ı,O���M&�X�%���^�Mıľ罝&�X�%�}�z��8���-�s��]u��\g3I��%�b{�צ�q,Kľ罝&�X�%�}�{:Mı,����>Oc�l ��?g���Mĳ��L���o�}]s���vU�_LK��=��7ı,E����&�X�%���^�Mı,K���i7�L�g|s�<��n8��F������v��1��s�x�%��	f��Ƽ$k�$Sn{��Jg8Γq,Kľ���&�X�%���^�Mı,K���h?O�b%�b~����n%�bX��lɌ���P��-�/�&q3��^�����ı,O{�٤�Kı=�{zMı,K���t���� �D�����ɉ0`�.1��A?{ߴhI�;�{��D����t��bX�'�s�q|q3��L���k��Q����2i7ı,Os�ޓq,Kľ�}�&�X�%��w^�Mı,�=���8�8���&qwwĐ$���V[&.3��Kı/��gI��%�b{�צ�q,K��=�Mı,K�﷤�Kı5����`�I��0w��JR���:wl�+� F����i��Wn�[l��g\=B$������𛲤
�Z,=�A<��R����lA�q$���r�H'�qڕ�h� N×t�%s�z�]�]\Q��Ȝ�e0m�m������cq���왉"ݓ`M�9;\�m� w/[��]I�<GT$��ۍ�SA�Ҋ�B8�B�1`ۇ�.A��*�+jl,��Y�n�&���A1�UB��T	\B�8"TK�����뱌�v@�u�{��w���|���M}��oq��K��^�Mı,K���i7ı,K�w��n%�bX������K�L���{��Z����L���g�b{���&�X�%�}�{:Mı,K���t��bX�'��zi7,K�������s��ۛ�d�n%�bX������Kı/��gI��?��"b'�{_��q,K�����M�&q3��]��qz�@㈩��s�ㅉg�(b&?~��:Mı,K����I��%�b{�צ�q,Kľ�s�㉜L�g��V�D�@f1��7ı,Ow���n%�bX����I��%�b_s�Γq,Kľ��s�㉜L�g��(zGGd�{.��^��{m�i�mck=ˮ�t��.JH0}ˊLu���ҧUL,������&qX�����Kı/��gI��%�b_{�Γq,K��{�M&�X�#8���5�T�;y-�q|q3��V%�=��7�!�9���%����7ı,Os���n%�bX����\_L�g8�����>u��[+��Mı,K���t��bX�'��zi7���1�~٤�Kı/��\���g8�ūw��B��Q�c��t��bY� �������Mı,K�}�f�q,Kľ罝&�X�%�}��:Mı,K�:O8�󛛜b�̸�f�q,K��;�Mı,K�)S���t�D�,K��gI��%�b{�צ�q,K��$����i�M�;u�h��KI�����9�:^�oN=����u���G��g3I��%�b_s�Γq,Kľ�}�&�X�%���^�Mı,K��x�/�&q3��]��qOJ&������I��%�b_s�ΓqTKı=���I��%�b{�צ�q,K�?w޹����&q3��w�++���$�g9Γq,K��{�M&�X�%���^�Mı��U�(�" ���ZEA���*�AdQr�B	`)�T%@�F�����HhP���������t��bX�%�{�:Mı��/��ͯ&WK`�m��/�&p��1����4��bX�%��߳��Kı/��gI��%�b{�צ�s��L�g���T��Go#���/�%�b_s�Γq,K��P��߿gI�Kı?{��4��bX�'��zi7ı,H��䷸�0z�rTir��β{t�ӝ�MƮ���0#i#n:�vz6����r�K��b�������bX������Kı=���I��%�b{�צ� Mı,K���t�L�g8�n���X㶊X�nۜ[�bX�'��zi7ı,O{���n%�bX������Kı/��gI������8�W���>������i7ı,O߿k��n%�bX������K,K���t��bX�'��l�n%�bX���[�y����9͹��f�q,K��9�cI��%�b_{�Γq,K��{�Mı,	�m���G��`f�A�O߿k��l�g8������=l㈩�-y��%�b_{�Γq,K���Mı,K���4��bX�'y�z�78���&q{J=��В���pŐ�]�ݶ0n�CK;�لۗ==�6.x��n�:�dN�Inq|q3��L���,Ḗ%�b{�צ�q,K��3�]�X�%�}�{:Mı,K�z��!���:�;m3�㉜L�g��zi7ı,N�>��n%�bX������Kı9���I�ؖ%�������ț����g�8���-�}��Kı/��gI��%�bs�צ�q,K����M&�X�%��o�	'�����㉜L��~���t��bX�'{_��q,K����M&�X�*؝�}��Kħ��?}v�Km�s�㉜L�q9���I��%�b{�צ�q,K��3�]&�X�%�}�{:Mı,K'|����	 �π�� 8�h����F� iYh���aH�+"� �h@�l l���|aʟ!��d�#+*��QC�q�\@�$�HF
X � ��BG�V��,��!�v�N�e 2d����kwhi���PJ;xs�i���D�\�{�j8	p�.g8�����V��P��[V점�m6�  8�7��h���Q! �zɶŶڲ�BMd��Z��X�/1�T����Ϋ����dCYg3�vK�K�E� �n��c�"Bu�y)rZz� B��������z��k��@jڌt�٭lڗ�*�pY�ݣ]Vvx|�b���8�%��0c5&�����u��mN�v�>�B��ggt��ŏ:q�q64����#C�v�ru���T����x'���fs��2�P��:�F�s[kk)Y�ծ[�M�ҡ��2WC�R�F�z�[
����<�T�U][U]FtncF��ܫ���L-�.��͆� m��v�s�.�%Z�u�p6�6 �)�v�x.�W��͍��ѵ�$�m�2�Q��n&�:�6��\���ql���U���
��H� �ت��"��p��Й9��M��)p6�;f����m��Bx�zĊӌZGu��!�>���56ܫ�u�[���:�!퀰�qq���e�}m���$�.��3�d��(�]���� Ftm����<�;[�F�����n��t�L瞐y|v�b���:E�^����0՞���&0&P��y2�fI�-��"ḅJ�Pbt�ֹĎ����$[{i��Ymݬ�`B��	P8��H6wB���S�����]��!�
�*.lc�p�mݷ3�Q��M0{[)#�b
�IFMٜB���w+u"�:�4���V��]�V�ۀ����z�խ��M�vVg�@�R��Ֆ,c��q�Ӆ�7XK.H Cu��V��NGؘ��W3��t���UI��L�λqe�Z�'Z�TsJ�[R�
�]%Ö��۳�e2@im����)����e�`���ѻR.�z%W�
X+��uT-Bޡ�n�i�0u�K�8-N�Զ�l�ݻf��U�h)i�\pGc�n�m�	�[U]�{�ղ������n�/sm�%�(s��q�1f3�ޡ����SnU�:tM���E6��� �#�o�:�`���T6�;����9$�c�F0;�W�v�u�iMx�m���Мh��6������5Q8V��c�]�Hu�Ĭ	�i%W6���U��Gf^;=�☠��Ը�<.�뤒2���q�]��5Xvu�x����<K���qien�yl���dzM),d�dΘ�ou����g����.8탗��YG�7`5�Ca:��(4���pj<���w���"���r!�qgFNZv���V�=�w9×���n�}��8wU��/$�J쪖Q�Oq~8���&q~�u��Kı;���I��%�b_{�΃�$A�&"X�'{��&�X�q3���o�O��R�ku�L���bX�'y�z�7ı,K�{��n%�bX��}�I��%�b{�צ�qQ�L�ggu������*j�^q|q8�%�}�{:Mı,K��4��bX�'��zi7ı,N�>��n%8���/��|����JF�Inq|qX�~ �������Mı,K����4��bX�'q�{Mı,�/��\���g8���{������:�c9�f�q,K����M&�X�%��羺Mı,K���t��bX�'woK��
HRB����{�����MU��\r�^��	ؖ��&51��Ӹ�,����71����}�ȭ�����7o#���/�8�K�Ͽ]&�X�%�}�{:Mı,K�{^�蘉bX��~���S8���-��9I%v�'e�-�8�ı,K�{��n;���� �l��K߻�M&�X�%���u��Kı;���I��bX�9�_l�d��)c��nq|q3��L���g���Kı=�k�I��%�bw�ﮓq,Kľ���&�X�%��N��1�K-�,�������&q3���x�/��,K��}t��bX�%����7İlO��zi7ı,Nx�-񏫑R�ku�L���g8�Żw�8��bX�����߳��%�bX���_��q,K����M&�X�%��V��x_8/�+h� ����x2�����]�8�n��O��.���7@2̘z,m����n��%�b_߿~Γq,K���צ�q,K����M&�X�%�����/�&q3��_���;KY�hs�t��bX�'��zi7ı,O{���n%�bX��{��Kı/��\��\g8�ų_���]-��8ɜ�&�X�%��{^�Mı,K��}t��c�'h"1�@`����"�` �0!T
A>��������Kı>�Mzi7ı,O�0{9�	s����&�q,K8�=���I��%�b_{�Γq,K��<k�I��%�����u\/�RB����O��9SU��1�3��&�X�%�}�{:Mı,K�xצ�q,K����M�f��L�vrzZ����Z��vVhָ�6Hבz��3�#���.ǷGj6-˿�����)c��o�~���n���;��������{� ��Q�e��,�,��сm�d��-�0/�*?���?-i�,��B�"t���w� 7wm���L�j�,��Vg�I�sD�W����XmՀ��2�m�V	%�%���_{�������@�'H��`_\T`[k��.�mL��~����)��2u���6�X��r7��׷<q��Wq&I�f�zYi�,۵`<�9�ۭ��75V����E�_#���U�ogu���a�{� ��+� ��ŞK�Cvy���؎MM*�U��{��X<T�=	L���,_w� ���=�X㶊X�n�Xj���zX����c�I(�������|���e���JIGU���j��I�z|��V�T�T$��&���r.]Z���[[ta]n��y�K��oa���p۵jΉ��'kݻ2=Bŏ]㨶�nzNƵ� ��<�N�:�h���X�U����5dWP3i�rNb�'M2��,۞8��H�v���*�H5�NzjN����g��NY�G��N;bw��=gs٣��ț�'mZ�v���Ïu��k(61��Zΰ��ۚkl�\��Z�8v!��x�v^�����z�s��}�U��d{n�fݒ"}� 2O�U����v�6CsR�F���V�NKm���|�����p�T���ݭ,�rOʩ�+�JP��S�qQ�mT`I~��uWH��Ѐ�-�>�WLwn�{������p�����^89,H`[UEFm�����{�<`^�5�E��t��{ۥ�6�XͧVn�`~K82D=͆�b�N'�CE�:z�=Z�q��������v��ڰ[�0=:��]:)��n�Հ|�u`6�I} ��ֵ�샮Kh������ۇ��r"&RHt��o� �u`gLC���KiK,r�pݺ`�n�{�\M���p���pں�z��NKm��$0$�u�[j`[�0-����X�֫g,
�,� n���s�O���~���w��`��0��mU��x nc��]N������ixܼ��瀔�h䭡Z#uʊ��VD�%�������0$���Si-�7��D�-V��t��q.$���\R��M�{��XͧVO(���rGo+���;��x��p�8��\�Ba>IA$hU�TJ��3�� ����׫ak���]V�l=
!$����XwVՀۦX��x�]i�A�%��:۶�۫nmT`M�� �������o�r�����[j�ql���;]���WfxNz�۶�`�Yi����s����1�h�R�X�V��֖Nc�6�XͧVZ�R�e��Wk���`��?/s�\�$�� wZڰ39�yBS'g�$�9U2$v�CW.`��&��Sڨ���v`~��Z:�dM:�In��?��B�s=��`{ޯOq��"a�"'�������PӮ��ȟ%��u�,��� m��>m;V��
#�v��ac����A��XÇ^�ok��Z���ŭ���օ!�[?�bM?�����F���Q��*h�� ��߹`��ӵ`<u� wWY5;lm�:�+�`�v�6���X9���"!)��9S�\��G]��p���,{�L��׀�ۀw��o2��\�$��U`<t�3���c����uo���/5�ZH�v��-����0sX<NՀ�ݫ興S�+�T��v`�;=4�5�|�U�J�&� ꣁ�w�;��SlN3Ǡ�{s��RF9�0�C�:Uܳhd��9xݧu��k�ة�D�#d��Z:��I;XvvK��c+;��{a������.�8�.ޭ�ݰZٗ����R��όR�N�e��N��a@J�&:��6nt�<e{x�i�öl��S�f�M��⪺.U���*������{�y/�V`2'"��綰^���D�؃��4�9��l\�ΥL�q�X⮌#+e��=��X<NՀ�ݯD(K�8��q���ȝ#C� �z���q`�� 7�۟�.6u�{�ۮ��dh�K����VNc�
#Д.p�������ŀj���N^H;y],� ��o0�S�r�`_J�K�J�J�3%)�\*j�`����Dy(����W@��Z�2s,9��a�**f��b�K�˧zϫ��Y}���J���z�3;C�����i�\��G[� ��]0��ŀu��0wn��o.��,�VJLL�jI߹��eD	 ��,8&�a���&ﹼ`}�������M���^�夊Wk��ʰ{�����%��o�� �wذ��Y!�W�\e`����n���`z~�}+��K��6�5]q:F�;n��.���ŀu��� ����ok�r'�$tvK69{t�[�����<�;=A���ע��֤������I��6�uYRRS����ŀ}:]`YS�AQ�3ֽ�Y��j_�P�c��� �ʘI��	�qg��a�Z�Q�a��dvW���gRM�{52at:G�ȇW�ғ<��7���+1A�T*�I�#uL a =#D��Q�RbY]d��5�S#�l�q5��r�,H:�LT3040Â����� O�N�>X�!Pr��v��u�����2��m�Ru  ���T�s��N���ԓ}�;u$�Z{��Imu�%� ��[� ���,���������=�=��9e��F��	�^0>�.������~���w��͠���`��F*E7j�R��[t��%��ϴc�Oc:�����(��p���P�g�z����*`}&W�K��/�=��ŀk�2C�т�eN��������^0'�x��t���ݺYZj��t��n�z����X{�M�پx���~f��6�u^qJ�R�V�J%�ߕ��ǳ`<u`y#���������8���1��4W)Xg1́�{�k�:��Vw, _��{ �6�mTv�ܵ_����6۞�x��n5Y���#�'ON�x����+�]Xiݺ�yaݫ���_Ɂ��^0/�x��������܍�Kh���-����_���羵`f�}6 ����7�h�:�%R�v�}��x&�w}p۫ذ[�ds+�����E��"��ٰǵ`}���v�~��t|+"��J�wm��
.�������>�c��� ��(��b$�*Ej��U0��}�$�Đ�s���{-ļQ+ĵ�=�(�⋌ۉ�bC�ۺ�� ���&��I��m����5����+=���)8 �ظ}�ca�j��r�
6n��OP� 	˰{1�)x��b3Oi�"dѳulzn:d�6�9F�t�Yڑv��S�2�q�n0S��h��H��@��ՠ��][N�۷YŇc'�.[2D���\n�Wt�L�r��'�IqU�����_1�����tg�!z�m۶����!0N�q�����X�f��V�c��V����#C,��~��V�S,����Q
>�7Ձ�i�Sn�Wi"�Z�X��� ����wn�z����8�������m,����q՛�z��V�0W��[��7S�;+��q�w}p[��0/���L��_n��r��S\�UU��bv�%��>�o� ��ۀo?��핢�v��\Yѐh��vt�s�nS�i����G<q�������d���+%�5*�7�n���� 7�v�/�~�^ŀy{��9��
Z�R��f���3٬���d9A"���rCq�XƶՀ����w8r��R2�9L ��ۀ}ޭŇ�8��v��?n�ߧu�[
��$�UXj�	%�f��X{^,�)���� ��5jm�J�$S��n}H��/�L�2�=0�z���n�q��=�p�[��n�Enw��Wl�^���6?���{�M���nx+��\��n���u`f'^ID%􇻾ŀ]������NTHݦ o�Jd:�ڰ7ڰ>̦_�$���Z����o$��-��uz���f�߁��
�Q���y(���eY`{�:����j��$�v$�����T`Ҧ��V j�Mꔰ���t�����l(S������`>�`z2�xO9��Q�3�;��6��;���;fE�Gh۴����N�[��e�.]k&��6��/���L��Q�=z*.[��8�#C,� �z�$�g������ ���3����3ɷlU�Q:�,`~�~�Q�w���2�`j���*��"v�[Ls���r{}��'��~Ƥ���Ԃ��RP#j4R#3��`<	 S��N.rOng� ���u�,q�9Q��q���Ifl���7i`gr�{o���|���I��s��6hָ���M�5�ʛ�6��Q�lEr�:)�.H�;����.Z���=?�0/��z*05����M��$����-d%X��x�������z�� �nm�du���$� ���0�w^����I);���,���X�~�$5��댯�^�Xz��zW�?�e����emV���,r���n,��5ﺺ��������@�(A  ��"6N�N���39$�gU�-�ȹ���Ӹv�&�7�r\hZ�Vvv���,;��ݽ���Z�\;U�0��Z��$p��-j�({\���	q�C�}?e�v�j�p�/g�6���N.�`urmn��W����J*r��ܻ�q����[s쁵��)1�vd�r$�$��h'e�i
�=R�$�p �a�9˕�b���NҼ�2� �Bk1H![�:}��������{����>� ��WiD�ܑ�x�݇I�<nW��b�q��W�����r=e�L5f����͏����	���l���ԯ=k�UJ��t�����\l�������Xwq`�ۮ��2�*$z���l���ЯҼ`}"�ܣ��,��-�ߺn,�����ۦ���=��|{�z�K+��i�,`OJ������ŀ}��<qV�q���":�=�s�۳���n��������s$�Ap�]],�9v�;�0>�Q���y���^~�����}� �;���U��]���y̝����W�	�^0'���EKK��q:F�;n��7��qa�o{�� {w� ���#�@��5<��X~Q;��+�,�:�z�1��,˻�qYybnZԐ����t`J����}k��SL?~ΰ�-);��R:�n�V��v��<��<���;��w��������dMpݔ*��{w�`w�.Հ�ݬ_Hw8����Q��Q�ۜ�W#���6�~�qXnS,�:�DD$�L�Usxp���j�S�U�{��,���\�g�9A `
���J%L���S'�C{�?{:�o��ѩ$��M�;J�l$� ���`��p�%ڰ���.y��V��	����ڷ�Z��0%Lzmx�������~���F��yS�m�\�'mmt�a�2�����3�۴��p�tkTdj;�,��MI0=���׌�Z`��p���$����')j�[�~�D%�8f�}6��U���X���qZ�brZԐ������%Lzmx���� ��un�\v�NЎKL%���7��\���������B3�ަ��t���嶸ݶ�o^��7��,m� 7�ۀwxD֣%���T�Gj���ewS�W'�pݙ�W� �T#�� N<�!m-�Yjqʰ��� ��t��u�IBJ;��l�Հyo�ϕR���X#�c��0%L���}�� ����sZ�2����0{ݸ�%ڳTBP����skK��2�l���41�p��q`�w������>g{�49-d��)+Kּ`_UFd����^0=����� 'Z
u*!LD)�"�H�A�U�X�Q~�� O����~�0�"S�"��UN#�����k�:T��B��& "�A2����4�>7;El�FY���B
�tT �hE��R0Xā�ʤ��5|�`K#�o�/o�����@8�ݔm�   p:Kk��%�[[I�D��Y/��m���43`*��mri6��	��LPq˶�c�}6s&͉�pK=Nj��n��c+�-�s���J�-��vz��D�\�q��ֽRq��2�.gc����ζ�%�I�j�,�������Md���]ڶNc�������[=B3���0�;l�r���M�:C�xCv�Z9����[��D�mGvM�:��$���B�X�7�.��ۋM[8��"
!��:C�=����m÷MA�G�O�[�Z�%���m�$�M�6�a��tmhN¢�+���%�m�� � [V��IFp��f�mY�]m��n�b�e���~��k��R�q��h[A�zM-t�<nuȱ�:sL���^t��l��7t�R��;s��tc�8��Y����m�?��=�Q�0횪A�n�#]s��l�$lr�l�'�R�2�Ŝ�6n����:�:��Opk�Ͷְ���"]g�`�ې�ݺ��;;j0�W63����R�9��%������x�G���a[n"�e��>'�t�J�g:�G�KԖ޵ۖ
R��vƝ�����%�"�(]��઺wgeU���ͮ��U��:NJr*� &������U���\�e8ZKn�\5u�	�v��� �m�͹ײ�:.Ƙ��i�'1uȉ(3�mU�Il0ݶ�d�R�u^t3n(�2\2mR�ԫA����nm$QTH�[p��n:U�a�[�o�������v@j����8�A[[n���xL;-�u�+gt��*J��P \M&s�nT�D��R�`�������/�p���
zڻGD�a�&Gm�6��
�\��`^�A�/\����vާ-/�)�G�m��te�6����6jͷ���-���C�[u'`�X�Ί�h
��+��YF�ݙO;��<Y:�LF�YkG6۔�mt �2)L�@S����  ?��@J�D���S�dW����x��<HeU:��vb���7"Yl��L��n^����hݳX:yk�oWt��.մ.L�m=`U��`HR���0@�l���Ƹ�I��3����n�3 ���3mçS��;��Ol9Ù��;�n��3��XrGF�֎q.�%���]�H��	�9I��nGV�n�U|��cl���z����)�n1��;'��צ��/V	b�S�����.-�&0\�ͷ��T ���I��eg�յ�W5��׶ݽ��Q���;�ubB�;�B��N4���\�߱�j���k�p������`J�Y���׌W��[���S�#�� 7�۟�$��;�vՁ��j�o��J���3����29�mq�m�;����`�w�Q	%3����k{V�dM>UQ�_˒����^0-���S�g��� o���v�mb���J��ڰ<�D�ݯ�������mY���w�/�a�	��rn���sz�՞�݉<]���\c\i^un�j#�N��[�[���S�v�`Yk����>�ۥR��$V��� �u�,�i�Q	�G�����s���@7��?��������"��Z�B���`kݵ`7�Հ<n���j�k��qZ�brZ�!mX_�\������o�V�˵`<nՀ5���Urd�ԃ�{�0-L�W�-x��ۦ sV�.�M��R�Z8;\u���/n����n�u+�����h���q[F׮��r1UU<��UX�;V��X��D~�{�����w���^Yk!*�7�~Q2n���5�Հ��j�d�>�ڝ����I*�=��, ���;���VJ�ap���E�E#+`��.��ڰ5�`uI��<sD�S�*xW)XjQ��{}�<�zՁe�������	ؖ-�I�U���j��%�~_��Հ<n�m�~��/;��ؚx9;Y���ɱ�6�z퇎��v��)v-��NH쁿�����J��U(S�*��kݵ`7�Հ<n�����5w��+T,d�H�-� ׎��L��ڰ74�V��X]m��l����*����7����߷�ŀ{��,�!c#����UXz%;�ߕ��vՀ�;VK��")���9�SBIr���>�{���9y]��� �׌ex�,�0/�^0>�����	�����jA�j��5�Q'�j��۹�H�C7bz���n+^kb�s�^0-L�W�-x����I6Q𬊸YV own{��l�|{���`��Y��?wo��mUdV"�I�U���ڰ7j�(��ݵ`��w�:�;,���')j�7����Q�Yj`_B�`\���K�Q�Y"���m� �O��_��t�,{�� �$��^.sf�ȵB@��[Ɏp땯]�&�l�F66l�s:٭��M�mb5�{#'&��뺙����;��:���$��Dp�:������N�1v�� n����m�n�ݪ�'n{vq�<5NI.���[�&�ە�p�=�F�9�q�ڕ��gԤ����V݃�Ĵ6��лl��+���U\p�I�v4�b:j�H�nQ�'q�m��ݺ��l?����}������sߕU�)A��4�۳�^�۶+��6����62nn�F��]rņ����"���o����Հ���`<n�(�]2��QֆO����r�\n�pwOb���M��{�������>��l�m-�Yk8�-x����	��`_B�`�������Д��m� ��|�pv�<�/(\�{�V���窧 Zv-弱�6���W�	mx��۸����ih�4�N��/Wn��yNͺ�&k�v�{�5pvn��R�ֹ��j�[�p��\���x��׌�^`{�0��V��岺�Br��	���5@�V�����O����y�z`����;����*Il!!m���`M�����[^0��trW`T�7%XK�g��{�?<`Kk���`}0��ۨ�q՛�s���[^0-��m���n��핅p�9#j�	EU#X�a6�:�[��t������ٺ�	�צSM�z��N�`cnՀ�ݫ%��/%�o��X�^�m�GiT%D��`�׌	��`_B�`Kk������k@VE\�U�u���7�Mņs���C) dT��P=�)�DJ6��PP������RO���ԇ���+j�b)Z$r����=��/�ߞ0/�x��m��.n�rZ�v����-�ּ`M���鸰�� �[,��,���H��å�I���q��8%�^+��vl�}���|=l(��8H[W�{��,�wf��n,��� 5~�trW`T�9%X�o0/�^0%���^0>�7�,p��J�ـo�7��Ň�9���{����;�w�2G\�Z*�IÔ�mڰ�j��m�¡%PD� I!	BJ$2��g�vw���]��Tv�BTJIV��ŀd��`>�ڰ1�j��BQ��s�x���n������=l��v���G��]lkm�y�rum�lZ�0���w��}
�Q�h�C������0/�^0%���^0>�t�-S�
�9f���Xww��ŀu���?~�V���X��J��ݫ�v��Q2�wy`ni���{��R[H[V��ŀd��`>�ڰ�K�ߕ�j�6�g�Wh�f��,`M�����[^07{�������z�m�-9%����q����..9ylf�7�v��N�D�Z��y֬��sB�/Jz��dQ�j��Ѯ�HlĪ�]�܅T1�r���)ĥ��qlA�yl�qc)ͧ ��e��g�pR�v�;vֲ��3LQg]ml�c��%���
�c!�Գ.�j�F[Us����ݯ���c9��I��E�r�&��{,u 79�$�2[3�~:�)��U��\��8�cHu�����Α6�cb�d�B�+n�3��d�c�-�n8�]E�.����0%���^0&�y����fH�KE]��� �����M���V�����j��DD)�ƞ��ҨUe$� ��ذ�ݘ��q`��X�~�M��P��YV�"!K������mX۵`c�j��w��mL�؅U	� ��7��%Ē{����mX-�X����ɞUtC�Cۂ�ɦۍ�{-�6-wE�V���'�=G��f�����&y{pڻ�m������5�0=�׽�NJ�l����ő.p�H�,H�:PR$�"�uc�����ڰ1�j�����8y?��R�N�������0�i��	mx�����Mͬ�F��i�Vv�����-��Q�6��t�nY!eN^Wk�J���,��9��ޟ �wy`w�]��Ls�s\�h!�C�=�N�ۏ&q�ݤX�v:���^;T.+J(�nUA�GiT��)%Xv�M��޻^0%������R\ ��f�䵁6��	&׌	mx����y��s���f��QX�B���Y�6�mX۵g�Ցj"�
RH��0��(�"��P(��oyӃ��~5�f!
�f�$kUB(�2���cH����!�B�"�wahA���*E���HP� @�{D��B�JX��� L"p�"C���p)�zw"��`�#B6�����pB �dV$��p�b�������i�|��0�:�c��b@�4�I��;�q��K�}����9�x��"��B�\��1$�lkT����$,�Y�!$a+���2f@��^
Q�|�d'D�DXh,H� �"8A�=@
䀧A��5��}��w����;c�8���V�{��;�ݛ%��R۝�X{�mB�Tr�BBڰ�M׀.%͛�πm�ڰ1�j��H�eR�Uv�����l�gm{�0۲D[��ru�L��X6n�S����S��k����32]��v�	}!����iʝ��F��Y�Wj�M�Z���ݰ���D(�I.p5x��&h�R�TT�ӹc����x��e��,�0$%x�;�Z*ݥV:���`>�� �n����!	d!!.yD)�B�Ñ�{�pԓ}��1{���T��ʮX����(�ǿ/�׻k ��v`�k�����"�m�%�I�rl�5�bD�0�9xx�x�E�D�mz�T4�m��B�� �N�,{�� ��v`�v����M��q�ԅ�X�~��P��'}�X�ޫ0�k?��.s�����mB��r�A�j�?;��0-L		^0,���
鼙\n�URWl���~�z����ݫ�	/B\��{�j�S�G+�2*Y�{�rL		^0,���� �v���p��%?/?/9Kkn��Y�ݦ�]\�{qc��q[N�c�T��c<C9ݷ
r�4���)
�k��b���ZȧU��E0�O;EU�c]gp� tvB0�3��f�u�]�֘�Q����.��m`��ը�<�����+�q��/�j}C�b�	��5��m@��#(Fn�6�),��O9��trg�8!�tv��ٵܹ�H�-�꯾\�p��>�r*&�R�l��#dC�_Svl�m�nԙ��n}�7J#��X3��>��*r�Y%_���ذ�wf ownޝ�X���qV�*u�%� �e����~��&���d��W�XB*��ـ�v������qq�n���0߻t%�6V۬����+���`}��a���?~L{kkɴ;c�8�q[V����>}�����钼`I7p���B����-lqո��۳\-ݭ�9���2�����D���*�G%nKW�~{�L ��0=2W�%x���.oƬ�2c��5$���θ��� =ʪdDBT����h���j��ݵ`}8�,�]i�#�6+U�7e���,{+��-�}j`)?�n�r����;�0,���� ��0=2W����qV��%� ��v`;�����V�v��6-���ʤ:��p(]�f7]6��ؓ�:��u�I�ugY�D��h�\KO����&�J�d��K�z*�v��57�`}���^0>�l���s�6og�^M��Ӱi��X�ڰ;�c�*���" P��T��_<�V؛�`}�;��*\���orX���]`֦��^07��Xw�aS�C��UP�W����<�{����}j��y�l0rn��ߵ�n���4j�/h�{/n��X|77��˫�N���m��pqY���dBi���׌%x���]`֦��ct��/,�RU�o{��ߧu��ݸߖ�,�M��[��WT��X����`֦��^0,�����k�YMY+���p�-�I';��Rut�#�Q�(! m���sx��RO��q�I��6V۬�n[�}�n��?��޿�������;�=�NC`ܣ�؛�w%��zۓa®۫�դ��9-���s:2�!��W�mX��M8�� ;�� ��w^ Kj`}���R����o%��$���]`ژ{-x��׏��_o��p���T%���޸ߖ�,?����X{7� �~]i�+i�J53\��>�nՀ�v�����fwwn ui�z7K*���U%X��,��9�۫��X\@BP�A����I'����TP�����}T�-Ծ{��{�cT�[����&p�Ŝkr�Y3p�z���ź���u�2��Ws��-��� �[�ݧv���8"brm,�^n�B�\Ʋ�gv�����Ky�M�:Aw^j=�D,=;��pN��z�b�|I!׌b��嵖܁p0�g<6
*h}إ�g=n��<lGG9�2[f�� �Kb�L�b�Ym��	�HV�Ij��^\ĳ���@~�2�e�nA�#���J)ٮ��k��[m�L�{��6���**:�DuIc�h�� �ݫ��z�CwvՀ��s�͚�Iسqw-`ژ{-x��׌{���&��}2�6V۬�n[�~���X۵g���s8�l��X||�i��r4�-Xww�Ӻ��ݸߴ�X��G��+
9+p�ڬ�1́�z����ڰ1�`z#��^���������Ef�ya��{"k��M���e�M77&�z80Ӱ�
���ɪ:������v�m��I/�ov��?3��Nz��9B���	��;�_�,�A �(UPD!$�I	r��ڰ]2�n����ݮT�唰�`����)�~�7wj��i��1��DҪ;V�.X��������̯n��?~�9��e�j�L ��� �̯Z�=۸N�0�Յ��M`x#]hۣ�c���Q ��q�hy�v��U�]=�A�����!,�_�o~���K^0'�� ��0=z�e�Ӓ��4ӵZ��w�Ӻ�������X��-�Vr�B�j�3��6��Y�%؈���(��)s�/ذ{}� ��ܪ'
���hB.Z�=mL���%��lW��?3W�s��ڊ�v[�}�[� �mx���u�zژ��o5�r��"g�9�]r:9��46ۓs�Lh��wl]��oj��wHqq$5K̍��N^YGT��7}���������^0	.P��m����`��ş�\l;�z���ذ�w��]��u�
�CUڰ���>x��6)��mXi`fk�G�+��I)[��{��I/�Jg�{�����XܦXT$�duDD5	s3fe�;��-M�%�i�j�`��`OEF�j`}fW��L*�z�����f��6�=nܶY+�o-�wc��q+cr!z��-��Nˊ��:��꫾;�� �n��'k��$����Z�7����*�+-G*��v���"d��ڰ3��^2F�T�Rm�ʬv;-�?{W�`�w���X��� ��y��IS��Z�R��I%-��Xڰ�ua�+ ���8��r�l� ���,�$�s��]����j���IB����*��T_� Uh "���T_� ��� U��+��TdP�AP�BBBP��P��B�T )P��B(��EBB	P�dBD	P��EB ��P�@T"EB*0 0DX��T"EB	P��T �aP�P�P�P��`1�@T"��T 
(Q"�P�@T ��b"�T �@T"�E�0P��bDT"@T DXP�$B DX�P�1DX�B+E��)E��B �Q�P��DX #P���*�@T"(1DX����`�Q �T � @T"1DX�DY d@����� *�� ��` EW� �� Uv��*�� U�� ��� U� "���_誠�������
�2��; ߸!^������y�?����	�� �
om 
  
 �H �� �   �p^�   �DR P(	��*T*�  ((*�%
    
P(B�Eϒ  !�w�P   
H3 ���������p{���b�����`����1��sg����|�
p$�n΋��׽���@uh[��A� |    �P(��|zd���k�A��R� ��d��#�� 0;6���ϼ a��ϜN>��H�����+[����2-��� ��@ P  8l�|�#v9^��G}��z@.�C�=2t��ӀI�d{�����_p
3����h����{�@=�}��'�� �>  
� � >�[��.� tr � � �� � 0 �w � d�AN�� ��@,� { i:K0 �A�)f �0 ` D f ރ�|J
 �6 ӟA��&��;�{����c��4�={�=8��r>� ���}���u��	��`��=��ӻ�:�        >�jzOT��RD�y4 110� 4�6�QR�      )��T�  ɠ     D�*�	�m) 4 �  0�j~�P�%*D� ` ��i��a��)$�!4�=!��$�G��d��S�C�����M0�_�2N���{���N��ʀ �A�_��` �#�DT?z
#�����EtB��/��� �$���:��\TA{����( �2q���~�������Z������     ��   ��5 �@�  ��� p�����wd  8-̈ �@�  ��2     � ��d 4 ���c
�1�a�$�� _�}T� } � "�@� K �� >��U�� Q�*�� ��� � �T>�	�U��@>��� P� D � /�TG� �@� �EW耠} >�
�@� ?@�
�qA~�� �lU~�
�E�� � �*��/�O��=@ � '�UO� �@<�����.���Iw��2���2�~+�ǭ>����/+�i4���3<%��G���f44��a�xy��q�3
��9�8@�hqVv�퀺 ��'a���w��|�|�}Ϲ��r�<�)���m�n�)×S0���bjP���\#.�C�DQ��B�*ե\6�,!��8�xK0��F�$ �K1]���<�#���$��4���WP�\��������ZNK�ә١�,*�=<��NoF���c�����I���$BD��Á�;�ip�aHP��H4#bH��:��Izﴄ� ��X2̅��
�3�'Y�8s	�M0�"e���jD��9�\48�z{cS8��9���#�a^��9�0��'2i��.��!B,!R"@ą��k7Is�v
����,L�^>7���Q\{\��]��0�+.u�k/����x�!��Q��#ST�F6Ǜ��T��t�Q���L�C�
Ċa � ��uޞy<�f�:;��o�
Z<��K�K�y�
ˈ�@O<=e2\�N=����2���O:���zFob;L�E�M�íA_{�=y��:ɮKM�HP�9�]y�w�4O8D
i�u��w�1(��R�b���)�2Ve�!����u��6s״"�"0���6)�X4=Zw��Ρ6�-H�
^���32C�xbPa 1#/gP�*\�Ji��F��N���|��s�y�L"��<)� v�&�^>.m�N�f�jh��P�aNzrxxe���%Ò@�
��/�q���t�s9�y$o]�5"Ab�4JB'-�K�),9���	N���C^#ڤ	k
�9;�64�Y�D*�= u^���b�"����H���I�C�鐕���Nu#$#�
`��"B$d199B2%�X�5�q�zcQ�H�i�jI���xO�c`RR!`�#Y������h��T9̓!\D�58��s�.ob�\ R4=<��WQ�P���Ǽ�YNi�79��	8�Isp�.;����F�D��8�L9���H��*M;�JA�.hB��w1��%L�B,,�$L�c �H�oGF!F5H/��)�3g}�7��;�� �ވz�=��!%�  �1|OX�<�$2n�g	{ó�n�8zz�A(`jq:NÏ�N��q���|��Ϊ`�;;z7zz����D��Sx$
�h���aN��g���F^����ކɭ� ����!X[X��0�P�i���BF�	�=�&��xh��#[k�z�Bht�Zf�H�/F��7�}`!�z�<Ğ��6�(��!o�u�}e�!�XHU%#	�ݡ9����E���ms�t��４w�����X�1mt��m!wt��ozs��Nv0�z�-D� D,�i��~t4��tB���� ^��Q�@"�a�M ���B<î�4E�GX�U4Yq�ǈF�F���GT�Pp1"T�T�
QpC�!�7&w�=�: �H6�p��CGML,Nͅrxi�Ǡ�C H\l��B�HD�X�*8��b�J�,h�"�+b��߃��w�!�5d�pz8�Ԟ��d"GHBI!'}�g}d1�Ι1B	SX��#�1��!E�;8z��C�Oo��z�0k��;κ�¥טr�`���Ì I"�k��8T�!H�RL��)��j�����k�`V73���;N�{	8�	��9�K�!��4%�M8p\��6�����ǔ{Π�`�j����H�`S$ׄ.!H�A�4�a��cE�Y �"D��R��HŁ��H�)B�(@%��2�T�P�e�qYR\%��HVP�M�CN v�� N��;à�@:y#;I!	 D��E�X쐬`�X��"D��=u�}�s�����M#B3;�:�{_A}띁$�z�c�8F)���B�%����i�!�u��N��a@#P�׸1� T�3N^�
�h51p)�0aq%��^�\h���,A��Q�ٮ����E�!J��.m��6gQ�\B� �d�(�1����d(@���+
���K�vn�C�߽dd�e����R6)p�3D��N�I�	C!�
L�0#:�Sc6�����i���wHҤMʛ�3X�7�]Z{�/G.� "���"U�RQ�dU0FL7{;6�|S!�%R-te뮎dC�:b%qӳ�;CS����W7z	�\��tM�#���C"@:�jp�y�n��0%1�LM�9���w��	�.��Ǟ���)
�햲L�Jl���*�0���aR]fic
�ƪhF�(HF�!��)�l17���i8i�˛��0�L7dQ�t��^@�:%��U:H�T�\'��o���FE��.i�J���o7}�%���H1�����ĀP�0��=�'~u�=<`Q#IV�!G @b���P�L"�x�7`2S	L D���H�LCF�KL��sL:
��Z��3N�~� q�1�Ț����i �Z��$)�$��i���K��!�{�:��N5W���B\�X�x� i�ID�4�*�^�u�F��4��Ilp�T00�B0�e�d�A
�
� @�$cJ�FD F'���Ӳ:Nt�	!iN���`L��*���)�6�!!��ŀ�`@=��$�(G�RV\4�8����݅�OEc �	^=��9����`gS�;��｝_p6C��5�6$ � �b@h�]V Q|���� z�>+P;�`g��R\f2�߭&rtޭ�V^�	�e�SKF1#���ā
°!�v�$*i�)�Y����#X0
w�4�o#�)�^����P8/L�CKK
X[��zb�5�4
 F�1u"�LCD�*��H5�py�ZK��#�*����ffݗa)�<n������.y�����L�����K/�=R��ӭ��:K����5k��y�v�-u��g�����<�ߌWo��&�|}<�p�}=��ִ�fl�s�0�~�����l���C�qҐ������YM6����z]zyε$�I$�I  H              �       $     �   �A�� ��� �  �� � m�  �  �  [@ ��         ��                                                                        !"Y]"�e�	vI�k�v<�m:�@�`Ѓ ���]�cv�j�S[p �%�Z6
N0lJ��W������\[e ��]-Xk*��]X1���Ά�!�F��ƾ��|Q2�!s���a���X*�ݺ,��p�FӋE�S���~[�-r��a�n�V�Ѫ��SS<�*Y�iI��R��o/<�Ll�6���%�56�����=��`�U�mP��j�  �2��p�ʆ�b�i`�ӯN�����[�l(�m��H�Հ   � `�+UJ�To;���LVͱS[��R��&N���! �l�������v����lA�T�'���_<�R�ݧjX+�pmv(@�e%ul&��$ -�l�Rf�b����@	 ���M'0[m� �Vܶ�p�ao���[��ɪٍrC׳�}��6�m�˭�      �@qm��8�e�H�$m�xж�p  ��{ﾽ�l 6�-�� ��U*յ�V�u֛Y�np-���ƺ\@��Vź��  q��D�@[m�2�l,��I0RJ6�6����� ��ж������-6 	m��*��S��fi����P[`�mm�  [\	  � �bN�\����d�F�l�A q G$��]n��im@appl�[@�v  -��[����`��dЎ�c]l�r��UT�	�̻S�6��ʺG���a��pI6�E��Ɗ�I���  �-��[m�[R�t�p��mmĎ   n�5���&:��[@m�� �W*� ���U��� BF6��[[ltm��aB��6lܛI���ܾi&����ʕ�$�c]Uҫ\�lHmp���J������]�n� ک\-�ړl�-l[@ i2�H�l8���[#$�e�����n@�"-6�4�*�����f�Uj���(
����y��R�]K�+T9iK7mml� �&5r�!�u���lT^!�LËo�rCn�Ͱrt    �&ҥ<��WUUK���YV�� o-n��scci5�\۞�<컲R��2�,<p[l�e�Kq��< S�ݧ����iY^�4�ܒ�t �J�W[U�mg=a�5�!@UB_6[nh4�L� �SIM�( �ܑ�ͳl� �0�   m� \�6�zඁ�cb���a��&�i���AA��yۥZ�����l*�Smͱ�k� ��IT��҅-ㆬ�'m<��YR� m�t��,�^�j��h��8&�/]���[m�h)K^[�l�-�&� �mC��m$x��)M)vH[@�mmJ����VҼ����]WA�r�V� ,u�Tm�^�8  � m��P V�K��ku� �4�;m�m�  [@��NH ��mYƷ�B�㐝8�@���m� 6�G-�|�v��l�H-�z�K5��v��'���Z՗��Ϸ�}��y%�$aH  �` 6�u�Y{u�m����.B�hluΞ�Eq]lv�5�ɵ�٢L�-�m��   �Xn�[�$s���кi1�lH��I�X$�#$C� � �nl�Ai�夒� pl� m�	&�8mx �
gm�vmP:%Z� �`     5���h8�ݫ�� ��p��� l���+i6�  9t��jtHM��m :�Jh�a����RPTɵ@H�n�kqn���[I ��q �p 8�Mk[Kh4PH���ä^9�zX�i��Ā�g�� �Îi���`8�u�p�Z �$I�T��%�\�� 8Hm��`iR�m	,���KoC8���I O����N�++U+�5J�ҭU�K��n��-�nI0��
����yYP �gj��v��s`$  4��^�jVV�� %��l0m�uK����8��We���Ϟ�^��-T��<�����9J����H�� x��n��K�Ͷ�� ��z�i�ګkh .U�nYWG���HꪩP�#\/Rm5�h	�Ekd&���p�"�G]`�_/�):��q��Ύ��877S�Β��y��n{+f�Fsk�ɲ��:��`	MИ-�Y� �OUV� mA���eRI �$�vy$۝�7&m��$��q#�lհ	� �� ��[�[ �%�젍�.�UP�����@ ��ﾸ�������n�Q�dm�(   շ� �-�� ��f�6��`�(�vN� ඖ�X`q' y ,ky�h�Ŵm� �   �@���h    @  6݁mk l @ m�D$kh��i)\6�9!���m����:[@	��k�  ��I��� �ڐ� k�մ[Cm� �i ��    �oQ�J-���~'�=���취  H��` -�8N ��Ŵ���E��  �4a'�L�ʹ�   � H    �vݴ�     �`�����nݸsm&� �   mm���z���`D� �  h        i �  �I�  ���[���is��;���{�m���"�FJH�]z�u��i1$�  8�8���   ����'���K�f��ӧ-�:6��.�[A�	 :�zԂCe��rl�� �	���]��VT21õ٭��[��VF�ZH�[%𐤝E�^�6��DG��]"�p�  ��  �ֻ�l�˵�  -���   [@ ۱�Ԓf�'lٴ���-��.�fm�	�� m�`  m���+�P���������?�(�N��-b��]Υ[xl  5�m� ��M�L�&H�h�t�H��]f��6�x�v� RN�i x 	:�6ٶ��$lV�[����U�U*Ȧ嶕'��m(�N�񰁰qJ����W[d���2@�֛lu	bݛl ���;�d��v��Ӏ.ڶ  45H6��N�[r�T]Pd�C�-$ZbHmȓ��n�Iv�h�ƻ:��P.�j���!̫���T�m U����r�    6�9m��l-�	 k�i1� �8[Cl��ؐ  m�  �m����s��k��l  ��EF�X��� Ce�	���x��<,e�2U� �d��cgC��\�T�s(�j�9�j��P-���mc�F�c������`�hi� pV� ��PF�l�먆��e�3,��7�����
(?����5Doh ��޲(�?���~ZY
Q$@�BBi��  �i�I��ci�L ZK��N��� XV������R R��))J4a�
?���!B�!B� B�!B�!  �@                       $�4$�HH	! '�O��N�T��������W�P=T�"�
,D��X��� �` c��8�
<F��Ҩ��Pb�b�c��y��ΐ5Q���uP<�OA|�uy�(�"<=<P
P�zG��@< SD����D� x���A�"z���EV$������
�b`C��:��\M�U�����CA"���r��\z�����">�C�"��{D;M�P�|�B�*�����=�)�:H*P<W��OAN����r	}C�L����!�p3�E�+� ��<LTA
��8 
"��LA{�(�x\H:��(� ���z	J�T��,=*�u�}$�@  @    !                                     ���ZI,%���0��I.c��ߏ7�o�fIP�{����y;-:�t����H��Q`(�B��H�`�E@��U*U`��fdφ����}?.�{}=[�\�ͭ�{�;�>��ߏd     [\� ��'��[Cm�            ��bE�JL��[.,r���N�/2�9�}sՒF{d�Zk�-�i*;!�ʱ[nŭ�;��ؗ�S���@mu�[�<�v��U&��"c��<�4�ݜK�L�s�pӒ�څ�U*�[��:���9%�S�ؠM��ڣ�(�� ��=��2�F���gWgz�9�&�9he�UU���S<T��؄UNة�,Ԩ	Gd4�-��ζH�2�nӲ:�(�[���-�ȇfݱ��9ڪ��힋�M 6�����t����K��{)H�d8V�Y`
8�We.�֧5�gdL��*�l�P������'e�4UW:3Ȝ�x�L��B���\�GKn���E[��tt�j�ms=��cz���fzn�Ɏ��p�UUV6;�a�4�t;5	�=�x�����{v���%e[�؍������d\�W��h����p�#����FҲ���7n���/\���+m�����z��]Z�Rc�Li�����cN�����ڝuUm'dح�
��؂��:�[U!+U[ud�Gm��>g#R�"vy�:�[{���)��R�C(U*հR� ��ee&6�ڕ`*�b��R��kwX���4���Z8����ݺ��I���c \�qv��N�6p�N�YS6�p��MVH�bEENF�)7Z�9t;[<�:�ۡ��v�y�R7@0�rĥFRt�`�Q�x�!��IUQ0�I��(�*�bl۫�F:Б;;���pr��@���M���.tf�x"�|�Pz�����zE�C�����x?  x��4�Mg|.���wsr�kX  Y׆�tP�%�k��W$�b�If�ئ M�����m�k6.kK�NtW�j۵���F�MN"v}ؤD��B;���q��;pt6�9�J�݊.�[���v���3��#)�3�[[�,����rGGG玸��M������wn⏝�w$�v�3���	.Jl���hN�0���s�д��e��O���j�[5�����3��&�:ж�we0�L����f^��<�3�=��+A�Մ���zk;��f�jd�$�`��E����X�E�2k�>�b:.�F�)]���st1��l����R���n�E�ۭӮ:�=�sA����q�s)�E+a	�=]�Q�4L	��ˆ�s̞wcLѶ�B�L�3xu��zQ�:Ht}1H�CõO==�k��Eηv�$i���5���;#� r{�v^��I�AmYe�l�s���n�̸i�f��xcA�����e6su��P��ic�����hW��q�NN]!���c�����s��N�m�H���2�8�n�v��;/M>�c����n�&#����,$�s&�����n�̸k���V��F�e�����`w7_ER�]RY/Md��A��ݻ`���n�̸i�5�wc�7e�PJ�	��e�܌s����0Ġv�`i��7|vM�9v�9zi9�2������4��h�Y{w�ȹ"$�����1����{X�X���se�����	O���Mw7X���sX��m�m�e��L�su�e�O��s�����m�N݆��̽4���wT#�0�PJ��T��C�߷N��'�dˡ�����d�dP�su���^�*�ve���۲/�k��&�ذ�
v��˷�u�k���\��=lZaI�]ݮ��y���3�E�2-��1J�Dn���s"����E�����ֶ��0�I�L�"dls2�\�d[�waJ�P��o��o���9�w���i+j�l��su���~}����z��>E��%Ip����FTC L�`��@t����`�q2�5S *1P(	����T��j�D�����۹l  ��,tz��XB�l�ƺ6�ua�r��i���v��q;Ʃ���ӃqbMs�@"�Ggm�]��7)H� f���S��u\� �nt��:9��n�*�V2ɱ�j��ul��[t�ANa�3�Vw6OX�\�b����"W�훦"44s9�]zc�e<�+��p!�vM��ⳛn����-�kht0�cV�2%��]n��5�.�r%�QUI)f[����>s&����3=�I���)��,$�rMc�����c�p�3���L����X�5���=��w.�Mc��@�%f�6
L���s&E�]ķ���n���Ӎ��P� �h��R�VMٺ*�\^H�u),<���/��oNv��2���Ю������I�ڶk�y��<��+ˍ�<��\5�9{Jŵi�d������c��i�k����m�e��n��U����5;�E�z�30+����-�
�I��k{KX��0�M�
kv.�e�:D6Vs���c��f��F�aɛ���-��/X��I���@s�1�l]�L'v�&j����c�������dv]�Bdݦ��fn�̸B��B;���l`Mͽ����m|/M<��3c���;�r�n���nٮI��dVk��qw��w-�w���M鱩+q�v�5a�]�3x<�\��S���Zv��پ�����.��s.y��m�*5m�l�XV��-=n�5�����1	5��o6�I*4�i7���@y��{5����F"��l��5�5�Ɏ�n��UP����(Q`T�r�m&k�ܳl]���v-5&�9ۆ�7�р޺,j��s�N6�m��96<�Y�4��m������8�d��\A�f���;p�f��P�7L�n�J�VѶx;��¨���Mn��Mc�I�c��t�[�m����Rlc�#M�s�gN^�Z%�M�e����$��{p�f��͸Jm[m�!�Zi�&�;ۀ�f����`pV�V���a�V]ݶ  �Zqw.���^k��\v��is�������jJ9��`��*�t�ƀ��d�5p�jo=�u�Wks��L6�i�C�ֳ�ݲ�f��ht����N�]�|�<�wl'F�\�]�c4��謎�]��[�U��ɺ��gkj���I�X��S���QeHY�n]�/�v>�x�����w�@�Tg���=�����nK�HA�m\M���ZM���3��lbf#VS6Z)��c�lc��k�;�l�i&�D��ݚ��c��Y���9�����6�&��n��c���ɣuh$���o��zk� l�聆$�c�0��b�W��Q4�v�Ui���]���ʌ��ZNa�84��Wm�m�5&�9/%ԛ7� ��ka2�A)ԑ���9��iq	$Z�@��(� ��PÛ��2��ɓ�m�V�m�l�ZM�n�xs.�c�%��I�M���e����^�̘�75&�'q���	��Lԛ�.���{|�Ȫx�L;�zI��ܹ���iq��a�� ���Ӧ�rGj��\H�ߎ������n��c�6$7d�vL	6?B��zjO�= `rzE�	�[f�e�ɏy�o�����\�8���}����߿t��+CzH@��4qBY���2BS_T0� ~EC�Ā��(��qS�1@�H�j��N���$� : A� Fb� 1�"B���c0!F0#E���s^���� ���b���IH�t���8%�J�r�N
wTmeUgp#��=RP�7��R!�?�@�����$ F+���(��艉UZ����! H!��g���@4���U�~P�+� Ρ�>�������C{�ǙU$UY̨զ_w�-�E~����d;��H��6�~
 �>���0$�c;p�f�c�  �.ֆHf�a�h��rG��գ{%��P��em��y��q�l�Mn���Y|�J����|�|�%z��I�.�j۷�����̌x�����o��j�0e����k썚���e���S���UPT��s"�W�ȹo���=�P���"Da�?>u�q�����:Lݧb�u��}��	5x�O�f��K}9��r�T�5�ܔ�X���2�y������$P��� G�(��R�����5���[�/¼=�]�0!QʑS�5������`N�1̹.��n��-Zm�����.%�Ⱥ�q��ȷu��S2IM0�L��s.�я̟{�}�'���9Q��']��n5��[�.�\;"�H�N�}|�����"��-浶�  ��sh픥f^��-tz�����f:y��O8Q�'	�#&{E�����c�`�+�lODI�ӎn3�u�Ld�i��;=�(�9�l��ȵ�smq����1����3��}���s]�^M�1jB���3#VJ�=S�ص=;9$�k
#�mU�pPm���Q��;��w���l����I��v�L�$yݼ��ݳغ5�\I���f nӵjŦl�S5��~1����~�9�3���F�M6�S��n�2l���LU��g����6��i��ь��]��9��7BeRA;)����]Ɍs602lc2�BYe�a���k&�9�02lc;p���H+P0]�L���G��ݶ6��\]�U��V{6+������M���k�7�`d�e��  ����\'Ki�wn݆�`d�o?@��~5��n�;ۉ{���G	RI��W���\����X�Q~�77ZV�I�-&�g3юvFM�s.�ܳ�I��)�w7X61Ò빸t�5Z`���$[���^�)�r�svp3GN��:�]���y���HN�+��M��=7,x�X�;�׎f�y�B	�O��{묛�}Y�����
�I�P��y�|����ֵ� A�R���>�r�t��Mi�t���O��}�p��{����we0�l�M�~U����@	�os��[K\��J�@�)��E��s���ۓb.��iɂ�:Y4�7&����Q���'��|�ɳ��妤�bvF�JӦZM+wRl~��ծ���y�;/�B���,�6�i6D�ތ�^5��z 隕I��;y�XH��*�B�dh� ��X�u��N�����e4W�|}���:����L�A"�m��:f�z������jOF�v�G"�T���=�ފ���P;�[��{1qGh����i!c���.�	�t�2�׽����� ��{�f�f����i�M���s����1Ò�3q�����we:m�$E��)��E����S�3NTm&�!���&�9�G[�/���zyyZ���[M��ԟO�> �� ���8a���/;���m��M�� *�����k�^+��\����E�[+4��4��{;�w4)�f�<#Ў�A��`_5v��'uڭĆ�WR�k�rl�4���s8ۖ+E�n�`N[4;��j�9�J�b�Ҝ..�ݮ&�����r�8YM�[�Ǟvⵛ�ZV�K.P�sǽ��w�����#��-���6�D��S^T8�gyy�ӽ�c�';\�C�8��sU*�%L^�ߦ�f{"�yp�=�sȰ�Dӻi�'��@U/��qs�K�9ϰ�#t��B��0﮽B��o8su'�"�iv�M;
�-��������cS�vBu�ݦݢ\ڀ̘Ǧ/�ю�-��ѳ��W$G���ٛ�vz����f�u�]���_V���Mݔ�V����̸k3�~��^�1����*��\����ޖ���,Z�`6�H� tr�c��5��f�V�$��E3�7}�f����/�Y:pDm��l�J|ڀ̘�v��f����"K	ݴ��g����=�yu��x�P���c�U
�j��d��nNڲ�n��E �r��n�E-�'�L��>w�;}����o��ϱ���Kv�M;
�v�I��UP� ��OO�;/��?Bu�ݦݣf����1��$�EP��|��*�7���=Z�B�f�`��n�kˆ�=���V��f�V]��m�{5xԛ��D4��c�E���a��V�qW9�8�0P�GD��=�W;4�Jc�+.�Ԛ)�ڪ��Vn��zpv_���,�,6�e�S�L�Y��ޚ��~9�<�0�,'m6�F﵉��i����@s�����-�S�AؼjM���i�P(q"E"���A�iRb�,"���yￛ�[�Ỏnm2�;f���$_'���j���g��q���7<q�	p�ێ�Ue�&�f�w+@��Dpj��Sv�v�-r�ګ�1�v/��7��}Z�V�SZU'����Rlu܊�����j�h[M�|fߍI��sʳ=�nE
F�tջl�|Fﵒ2j���K�d���i6Z ��Y<���pd�x�/�{5�o|:�vf9 @<]������T�s�$6B��{8����E����t�EF#�@�� E`��3Rb��U�bĈ(k��y		�䓉!'�لH�bC���D��I���b0 ��W+E�I��
�I�7�	�K�f��$7�����54`��HH0� ��E�0�X$H��b��d�	He��B�:�Xq�0�@ m+�
�q�Sf�Pb�Vܐ  � �	I!�V��oPp� �              z��V3Kr��}���d'*��`}��˽I�6��,#�բ��֎֎��۔㫶W�^h����-h��i�noB&�C/�6�Dsu����U[L�q��*��(#-P<t!;� {& b�I�pU��EU �j�����J.�v�Qv6��9���ؤ�0ܽ^�Z\l��"Z�v�"�p�k]
�M����YT�OZ��x����:B��ا��m+�a;ec�:�Vއ��y.l�����G�Ù�^پ�1�c�~������q�@��M�-\�����!j"�]������<���m��#�nUr�S��$��kTN�<��s�S��6�q�m�ZtQT�b�g�X��
�g�g�ͭ�WL�UU�lKرl�nܑEta0�b)�{��5t�����R䰅u�\����\[��\�I��!�K���l��U�����47gR�e�����8��<]���7`.gb�.i��Z�"kls�O ��B�WV�6���C5Y���֓�l�R� U@Rs@ �� ��s��Kn�/Zx��'X$��wK.��NU*tl�/3JKWj����l�Zm���6	S� :G��򖇴��/M�q�"&�m�˳f�#f��V�K�i�i�:�F]K+�K��G4�z7N�w`	�V�j��[`r���xݸ�hۅ�n�i�jr��$��N��ȼ��إh������Cm�(ʲ�I'32��-����q��1��J�#v�sv��q����� �wMU�A�W�u9���h$�_>�ȷ���{�m�  t�v��jn.%����w:ǚ�f+0�*�f�0�\����ᵞ���x�Պ�v�IS$t٧�Z6!�l�ӭ�2Ӽ)���g�u�Wqua�Bz�<d�X��Akg��&9�:-�R'�6&\E�yWh%V���t ]χ���xzC�
:�6ys&��Hn��n7fۛ�J�DZÆ��$.	�n{Rm�U7O;q�F�Tnx�m�=:����Gi�a%���*�~��ܽ5�zr�yW9�e�v�vȶ�O�K��H"M����`c	�x[TSw`�ڶjM�r��>@Q��"�"��{Iw�=
�ԑѴ������U���e�G��яi��M�I�J`�J��c�-5'��I�u�{�a�UZw<]mU�p���|��S� ��[����8�����+-�m6�=��Y��'�"OF=5��N��3Rz?�@D@���k3싽���н�y穲(��Ni��w&=2_Ʋz1��y�2K��	44Q���%�����@t��Vg�7RUeI�#������GXg��.��r
&��ܪU1��q���)��m�f��y�� ��KA�>�4�a%V�"�p>.���D��OO�h t�����2��۴l�\�>^�l|9/Ƥ��Z(Uϵz�r�N�^�ދ�v/�%ė�!j�W�B�=��[�*�����j�j����a^E�d�[��1\�dV]���e�6�e0iɌtV��b3c��L~{�~�^��PB�.܂�#]�nt����[�8�n������_,�I�Z%>�� �d�3���D*ON|{�o�0��4�i2����s.����Q��h4�i�m�m��$����Y��8*���IU�ȻM�#�w��7Uf{�Up(B��b��1����Uc �`�PI� 1��y���-	�M�F͵���U�6pv_�f{�~�<뭺�\]2�}¥	za�7����Z���ɜ:B�v�l��)��U�cˆ��1���V��/JH�)9$��[��yp���=�0�����;�l4�3��5 /2�w���l�Q���
�a����@;y�׈;��f��2N�I�rk���v� �}P�D���/�)�HޝF�b�  �mӅљS�k�nN:�Tv��S��4$�:;u�e݌0���.���[�l�D��Ԧ-�J�& ��q�z2B\���_���_�z��Cn;�ٗ��Wt��˞,	Y��1r�8��9]��)E	l��1E��Cb���U���f����{�{�����&m�.�Մ����mR,�Ջ���ܫL��PN��-<����>��@;ۊ[}�_ŭ�E33���ʪ�*D'tl���kH`]�@��}� ����|�¤u$t1�[ ��@;ۚ�w������n�!R6ʈ�U�6fz(�aش����W�y��E)"r4�IK`]׈��&�t�y<��]������h�o�;'lK���"rt��{c����k�g.:�Gk6b�b�UMF�T6g�P��͍��E ��v�-
A�#t�.�S� 0��`�2��,���2L���� U]��?h��;i�I5�N��2Ndj��(��@7�����#��R��� �� ;ܨ}��y�T��N�*&�'��A�v��E �+�wT�ը�ӨISS}�����g��U�
������c��G \��b�@9ۊ�Vw"�w;%H�@*k�$u�/=�Z�g;^ ������y��E)"jF䒖���v�?�oI.%�gި9�P�w�R�QB�*�m@���Ƞ~ִ�w]�{19�R��IT¢��*��P�c�s�����O3���Nw��k�Y��y 9벤[�ݯ�(��9�k��S�J�R����(_-�=��k`�ߕ�*�Tӥ�����64�y���T������N�*&�2Sߛ7y�n�����9��T����9K`yPv�u>��'�;\��Q��F�9���ٛ��aQ�|�g�@�� �} �}P���(�q�2�	Q7�M�&:�&�<[JIs��kLn��9�=Wƚ{����@7w �}P>w�o������u!N)P�܊�w��/���׈�i�B�'$)Ų�.����(|�TKR��L�Xd���ςh�`4�i:��E �� �\P�ʀq�$uD��"�E�-�8n�;YP�"�l����-$���[,~�I*������  ��v�rG��x.���(&z�h�*�N�
��"盞	L��;(�8s����념kK�Ҷ�cu������%�x�O�7� ������1��y�����Fj�5C��gm�;�sI��m���7f���Lss�Dm�gt�UwUK��� �1!�%��w�����u݌,۷��������3�qvų7q3���3�5�-p���1��;E ;ۨy�_Ͱ�׈,�2ERF��T���}Ƞ�x�w���M;�u*!��q�_��v�}q@w� �e�**UGK`v�n��T��w�m@=x��ES���
�[�ϕ}�v�dɞ��'�x�O�C�T#�j��V�%��-�"����{ѝ�d�i�ܱە�!���t�*��|�zT����x�l/�1O�Mi0�Mp�����1T �ׂ-O��ъ�W���������Q���L֒cv�+�KH���e1�L���;7x8~�J[K~��Ϣ�[ݧT�8��%:7�����v�(y�f�O�<@9g�JrR�#Tܪ���P<ŭj��[�^ �� �]���F5*C�3&;lh�8��ø��ޙř�tk�J�~����'X(��:I��'��{vg�����(u7�P���T$�*��%-�ۯ�n�s��ȧ�M�������
���l��4�Eq�k���3��}�}�{�ޏX�P��4%@�p.�>Ny�T2g�4MX�XH.� �p^�� F Bm����
ؤ�(��ĩ)�	�A�[�ˬ�9)�,	 %A��j'"/:���C��D4 ���yF "�  g���>)�� �����*��!�!�/��1���<S�Bt�i.�ۊ�^ �[e�PN�m9��Ϸ��}Ƞ�x�w�5 �+�D��B�R����"�o�� �k`v�����}���Cj�ʍ��Mk��g�m��V�c��]lO/��,75@�W��q@9ߠym�;ﶠλ�Q��IN��~Ƞ����E �k����=2S��I��j�"���w�[[6�}�� �dP{���JnF�M2�[���Y �\PG�-�Ϻ�?��H�H�T�n�.���v��Ƞ�E �*M��)T\b�,�pv�]���1�{	.�<�ԁ�t��
r��/2(;q@;�"���u���f�EU#iȶ}�P��s���3k`K컢S��UN.�oۢ۬ �� �}�gKd��:���E�;u��q@���j�寶���J�Q��7F���(���������(;^ �4�k�R��H�Z�DV�R b�V��!�o��swv�{x�m�  �/m9" ��k���y.iS�5����I���Hڌ��m��A�gc�Z���1��I� �Ls��6�;OdA������$ִ;��V�U�s���N�ѹ!Scd�t굃��4�;�i��we;\�d�n0�tY.�=p������8K��L���8!̻/4��1�{�.��cc��h˹�x<�]#��պ� 4��JI)Sr�t}�P��s���w��\��JrM:Q2�l֛��� �E{a۬&6y���P�T�D�c���I���T�E��3<���⺡�HAG!P��ͭ��x�|��ۯv�{�!�$�J�-��~p�s��1+�mm�WU����m��N� �tS���ϝ:St-�S76���JMԢS�P��MJ�`e׈;Woxٞ���[�q�+���RBQ�;u�sk���-%��l�v(;��6w�� ��J��&�Jtl̊��p�s��}2�*��$���T������do��=ا�;�ٸT�N�M�{@_k;V@;���nդ�u7-@�*:��Q�JB��<��<g�ۍH	�.�	�:�6�h��m�u�r�(;X@7���K�C����B��6_����@9u��׈{1��5U*U'Qp�� �*�~��/@�*����^�~M�s�����%9E
8JnC`_k���� �\P�q���u
UU	F����� �kyن��ǒ
;Pq<��M�6�8
(y��6���=�rj:z�h;�	T��
��F��Ƞ� �f>n�@9���T����<�ȸ�x�o��l�x�w���M�
�4TLtn6r�d{�X@=��{Sl;u� ix��	TII�*��;u���Pv�P>J������I%{��`{���U$z�B��.�(.�o��l]a Wm�n����q��R;>�����q���b�{Sg7 ^����������m�]�o`w+���E�ˬ��T���u)��|l���/+��q@9�E>I��yf��J��u!�/+��;wo����f���^o�*�!S�G�F{�����P��6N�x�r�͹U"�Q�m�[ב@=۽�ԓ�3�N��rl���$P���$Qj�QO<��s��Jn�ٶ�  ;I���Z:\�`j�Yɖ��n��	.�IJ-n,:M�	*l=�D��5��]R7��qIn����
�ث�s���v��"�Q��*��ecX�m�d�3���ͺ6��o�����{�=en
s��֩j�e�[۴H��٪�F������&�N��9Ƌ����H[�t�\�.��3e�.{cv�%�ۓ�q�ԭ�\�3�[��i�^�޸�g�O���kn�l��P<3P�D����������U�E �=����6�כg��HTh����E �ܢ��x���we�Snj��"��a���ڀv�a�9���k�-��'bߓI��;M$��'${��۸�����������T��WvN��Xx��Xc���zM���[�����������Du
U$N�,�|@3J�6�ֲ+��v�x������Q��IN��y�?�XVU
έa�rc��'��_�I6r�͹N��Q�m�[���`v�a�6_�	��̊�\��bu&��ӥ��i'y��;��۸�q�U^ͨ���J�JN9��׈4��� ��_m�n����yS�N0��}3xG �v���<��1��m���2X������]�%=���>�����M�x�f,ͦۚ�*H����J'��۫0�6fW��E<�w�yR�:��rSN���<l�a�f�������y�@;~�_)yK!B�I���;���y�@/���n�����~�)Tq��IN��y�@>�o6�m���k`^W� ���;�T�������g�2�9��zw8�٠��*����}���\�1�� ��Pw���7ۯ�� �vU�PZn�b�C���x9�P���|Y'=��� c���EBURrJ�l�� ��Y���}�E �߶���uEDIH�Hl=�$�����o"�s����?A���X@�R�=�����,�&ۚ�*H���q�TP>b����qp���n�q�g|�Aa�Gx�K�w9��$��^hz�6��CJ:�]����5Tt�RSq�Qp���������Kl;~Q@8זa��H�����P���0�9<�$�$�����z��"�Q��IN��3ފ��P�i��3k`^W�v�ܪ*:��ܥ�o�֓�}� �{�[�_>KO�{P��4��4*��Kdoי��/�����M�m�cORsž]��H��=�p,	E�a��>���1
D�AHA�D��4�U}^�=� ��M`��	x�rIXx�@	ЃR"��D,P)�XH��H@�¢�=
��xw<] �"���H��)�4�Ћ oI����/f ��X�F�"d=�'��C�jDdFT�U�!0��FR(�$�ot���&  cX�&������w����մ  l�)'V��Ëz� �              ����j������	�7:GL�,N����,We�s����pV��S�m�6���ۘJn赹�Hъ\�Y�cp��4شtlE�:n��
l�iV�ܲ�;+,S.��\Y�e�R�$fx*�af��t9����"]*��gli'��ld��.�.���A��%�[YE��jrr���hEL��Nl�)7m:�#a��7k�]�S��8C�� ]��8�iN������� s�v��5n�L-=n�یq�Xa��![���.�.����W"�Jʭ(��kF䘹��p���r,V���������"7��q��d���mȌ�A@Z�����P��,2��n,ɳ�#o� c"�Z�l�#���UQB�ٞ�
���6�'8�\�n�ָ��2skd��8ҥ՘x�&�2u����.܋˳g��md�kI�9��ԯe��Ix��ܵ�Yu��\F�Q*��E-������n��V{\��uu�í��^�ed�l�3lfW�A�,�J���P(��!��Ъ�U�*�Vw\P  !�l4v�egZ��
nR[�0$M�����4[� D�c=���� �ZS%�T�*ҭUUVQ�VT���&ɢu��rQղ��U;�"���mpnÝ[T��"��H
F�n]֣uH-�܊���*�ʫ!2c��1vd�C�>��dXPˡu=�������b8�	�족\��Ԇk1«�NsS�(q�u��N��$U��nffr\�f哝�������Zz���� ~��8�@����P⇝ b�
��hD����Y��_7v�2m�b�  �6���Mk �\����d�yPJ%m�4i�Xә."�tH�G;%ֆ��6i�d��.{��n)q����c���;v���Omj�N.ȆM��ɗ�ֻb���fu-��=�]g8���bev�"�,R�Ut����D8*ڶj-[�����k�}����b6yD���<�7=�;Eϓ�.[rY��ۛ��׽�����y���,�^ �b�7��-���fml�~�y�t�B������ml�E �n��n�@;�ح�朕$T�/q�碀e�ml�x�s���Wr�Q(�F���-��������+�v�(�~ڀq�,��)I UE�;u��n���E �n�����H`�T�����l�#��Ҧ�h����+���gG�|�c�b�&գ�����܌2O�'���;;��d��x��֒v�h+�R\c���a����OE��*��X��{;�s:ߍ�^��;}�~l��:�T��Q2�l1���`v�n�s���T�*�ӒUCv�uXC��2(o�j������x�Γ��C���l̊Z\��l���۬'�1��y5)��͍i�xL���`:�9xv�;�َ�) �q! ^$�"��`^z(;�f��׏����"�}�3ꔪP���E�/2|l�a ��Pw"�m�Wd#�R�EU!�'~g�d������<~<�T����0�>�p�ؾ7�4H��V�^dPv�s��l�a �N�p��J���)l�M@>]���C�Ƞ�j#��T��Rj�$q&c�:�qu������ܕ�e�3��n2��o���~����8�u��ߢ�y�x���R�rJ�l�x�I��"�v������a�z���U��D��aﾊ�GhXY�v�m���ePdt*�M�J�*���}�}Ű/2x�����/j��NI�hQ�%��~�9'/���F�*mG%7Ql̟��۬ ۽��~��E �I$��ZXC_@Q�,��ی;EˡW��8r\�-�mt^%~��������)$UR=_�� �~���a�6ui,���%)%�Jtl���$�������T�'��������Z�۫v�h+�hp�7�?��H�𾊠))�� �dP{��)�NA9I�K`v�x���۸�y---&v���<�
�ҩM5$����@/2(;�I�}�ӒM�U��>�H2Ys>�nM۴�m�  ,]�Q;�Ȝ#ѧ�O*���c&U�wV�e��8ͨ��6��7g�Nӹ�w���N��t�Cgn�`�G���#�ջ\�ۇ���ۉw\X�[mWa뭽H�գ���RaX��]�U\�]��li�[&x��n�����]�˳#Ͱ��rf۷fI����"fi��j�cT^�j�5�ׄ�IM��ŧ�=�%;4��Dn j�t�U%��(;q@9�Ϗ� | �Ww�_I����L�M��[��S�-%����6�x�v�)�|����U����H1G%7Ql�����y^!kM�R�9�E �^]�AT�Q��KI>�� �d_m�o�������G�$jGj��F��Ƞ-kI.�ml���^ �]�pQ�Ws�v��h݀u<[.�N�=Xi�^��ƹ�%*R�ۆ���Pw�ͅ>��䴗�Z�\��V�!G�eI�&U-���O��J����$���z� \��;D头��xZ�P��F����^ y0��E �{<lו�ۥQTh�Hl<���O�E �{<n�E�x�]ՎӨ
��"����ml��V�8�@;ud���~�(�p��玹�Px,��ǔ1v�di[Y��t�m�/bX� T[�s�۬9������v���k�0�r*RH��6cw��~�g|�Y�U�O��,��������Fy�h6�A6�g���;�x8 ��|��wKk����`{���o�U��'�)Rm�m�'y��۹���׈-J�=��d(�Ԩ')T�g^d��Ҽ���q秅 �Ƞ�ܵ6�-k5�<���<=d�;�N$N���6�M��J*RRr4�P��� �՞�ߢ���� �z�Ct�U�C`^dS�$�}��"�v�x��^'�M�����9$R����>���y^ ���W��eHމ T[kI�f�-�y^ ���$���Z�(v�I�����yϷ�g����d$��J�UHly�f���ml�E �{<l��n
8Tb#UE&�N�c�(�uبk�Z��N�ڱ)h1v���s�F��̊ �wQ@9��׵�%��ǋ��,�����)Sr�`g��o����.z�'20�*���
��j>E�i�jM2�[:�{>������P��@;���))9r)R-����-<��M�'3�2~��/$�������( �Q�)#�u�R��/��֖g��w���ǟ8�_�4��	ujѯ{n����܍�  [z�E�^�nU�咭�f�\L���e.ݱ�^
a�J�l�h�<�/P�=)s4B�����l;E�+q.���A��k�3N�M"�K��Cl�����9y��`�&��*�۪ۑ,E�9M��U�so\ݵ݇��;r�����L�Ph�ݐ�ه�? �/@�t[�D��$S#,�g>s'ݜsiN��V����K����u���&����Qx}�@9�����x�-i$���"�uk��7U�IM���y�޶;�v�({觴���g�P��R�"���<��6�kIf}��;w�����}��P�Rq�S���������������-f㪎J���)l�E�������L�ȡ���~�M�j('R�T�Q΍��;S���Ժw��[b)��n�������??�����\�'��n�ζ;�������W���)9%T6<󟒽*�RQ B�PR!C�P��x�
��??4�'��l����g?E��=^
T�j�DRG����mlAw�Bִ�o�s�ly� �W��U5*-�w��eǳ���8-.$�z�� �����8�@��n����-iieg���Ƞ9��
9R�����g��X�0�e�'���V�B�2�v�������_)���"������q@;ߢ��>����r��"���:UT�3"�֓e�E�����1�}:���[n�
��$��'���+Et��}���� �P?4��o�I�&�Df>�xs
�0�p��:O�D1A�J�T=q�"BVVM����S6x���707�:L!GCI�#�aTr� q��N��D�~��?�!��O�o��)ee���̓$��[qa��	U@!�Ã��eB�L���
�CC���tB�:0���@�!L!L40�����@��
��B](�H�:��! B �Ū�P�N`�{)$���i,k+�T~�U�qF�\%pyqԩMT��K��]u*�{������q@;ߢ�z�b"��%'$�� ����ik���g Ͻ(�s��#`_�i?�lN��ݳ:軲*:wr�s{�Y��m�Q��$�EJ�@U H��E ��Pw�k\1ߜ6ݬa���*��������e�O���͗�ޖ�;ڿ�8S"D������`[�8��P�� �X�jG*(�H�T���I<��d���$���2�
ʠV 2�I뻭��`w��*�*�d��/2(n�s��l}� ���̪T�7�Q�����9�����U��4�iҞ͊7��w}�T�)T��{�V���}���l}��;w�]�t�P��UC��0���|ִ�cx��y�@;��R�DU(D����#`[�8y�̊KZZM߲(n獁��X�R�
F�=��I<�������?��Z�e_��;�XЭ�6�t�$�k��UUd���1ߜ�q@?/,֒��>:􍦏,[@  �d����l�Ҷ�auyN��d�)�ж�A3 ț&����/��Yjؓ��*��+���흓D�%��Hu�X�pm���z��I��ԘY#۞;^NȞu���Y]�p]���-:�bGi��D��'��3ԖKd�۬���ut]��ŎΛ�Z,�W~s��>�ڙm���
xNNy��9�Զ�|�BD�&�tu��{���_|�d�ݩ
qp}��l}� ��P�� �\��#�"�EU!�-��q|��}{��$����B�U@ ;�O���B����=��[�"�o�{�����U�-���*:j�r���Iii��m@;w0���Ͱ�Ƞ��[�J���'-�۹���5�--e_���Ƞ�� �ikלR�	�*uM���eܻ�^�
Zv�`�-�,�mld��#<ݮgjzhm�1ߜ�q@;��%�|�3�}�ʕ*��n)#��0����Z�ZĴ���KZһ*v(����ߜ<�fAzt��N�c��������� U&�ߜk;�[��e ���8�#��������p���Z֓�f� ��������!�-���a�=��z(�w��:cx��=QPU?�cΰ����Sl���\��guǐ�[L�&�4��3ފ۸�7���_kKK�1ߜ�g,���Iʍ�&۔��zx��3k`c�p]�=��l�U�'Pr���2����ml�x��wo��,���w�(��d����M���;UW�}l�̊~Ƞ5��w�����x*��)�H��E ��S������>ZK+��ɨ��RS ���ʩ�!�2v:�9O/�$���?
���ĭ:JէM1��}�����6�����y���e"�I�
ql̞7�&Ǖ~{�W��|��f5�#�G%B9T���8{g�J}�2O$~��'"'�KM�����/��q@7��6��Ok ���������O����9Q*2
��K�gr(�ir�xpw� �n(��]��Ǒ7(�Rf)�dqa�v:�qu��i�g�`玌����6�#��;�<l}� �+���-o\�Ͻ>)g�U($��J1�w�]����2O3� �����|,XT��B��}��Ao���6���}�5USR�2��H��"�o��l}��;�ڀw��:#Du"-�˹�`u�8n�s������֒ח�ߦ�R��uֶ�  z���h�����t��-��Z�-J�U��҆$N�0���Ӳ�s�#.�SW��-E�7l�y���<�n�6*1�e�k<��Y��q]qm��%vf�=h&���:-$ٴ�d�u%.}kAr�c��v) �P��-WZ�UZ��3}���[���]����ݧ���x���l\��:���;>Xͥ5�S�;���o��I:M҅���:�;ۊ�zQϗ{�6^R=��R�Lj2S�#=��� �{<l��<���/ʪ"��R����/=5 �{,��Zn�|��>n��r9*	�A9Ka��U��>6?|�M��(����R�C��UIT��w��W�Ƞ�f�Ro3QBT���PU:�#h��+c���9:y���Mv��TQ���������R�q����3ފ��|��:����X�jUS����U�^��ib��֒��'����8;q@9����4GRht�;s���y������P��@6��jG%B:�ozIk_i$�'�p�����(���9�C���B�����=��>���4��y�.���cv�� �5��~ �
��Rhi�p��F�#g�Nu{���.�G��8u+�#�U����>���f���>{�"�ý��N�*A:���;۞7奭i��y�.�(������bdr�r�T8���'�y�����+@/̉�~�W�(W�|?*�
��x�'>���'�u�)�ӌ�H�fE 9ۨww��y�NLp�I�IZt�$��'�B��a$�@j��wW�B��m�b�ŵ���뀲.C��cO6}��H(n��`��y9��撐�qԀ�p]�k`[�p���I%�����ol8�|�u*S�C`c�9m��( �}��o䖓go"=A$��uT�Nm���}�-kKZI���y�7glܪ���*�-�kZZy�ڀ]��`[�8��>��D��E��W��|��d�S�J�N�������]�S͗~�~X���#N���m���n켘�S��=a)Hz�\�N�{luv#D�D���y�32({�-ikl.�x��OR)M8Ȥ�~l~���w�2L��e�[� �3c�i'M"R�r-����e�1�y� �Ƞ�g�!�m8�H��6�I�f�6�W�{3"��f���3�(����#�R���P��� ��P<�����獍�D�*o�%w�"� 
����,5[J�ґ$bB��JFƅ :D��i!꽝-�(�I Hq4 �L
�XzF�$X��a[�h��:/n$LDq)E�\@$[� X�HE�@��vpP�8X�TP��;��.yg��ar��v�wo5�Ӧ{m    8mrD��$8���!� -�              q\��ZUk�[�ב����GTu;''���Ϋ�8e���F��"U
۟7[*\�Uj��t�՛K�،��]��yz��1n�pl�k�ij��"�J�&�F�x!��`�����v�VVNڪƤ!�V�H��9r\Jx�&�e��e9sC�Nr�@pV5&^���6��5rlŪx�&�#�p�E�LD����o(�wh��0r��Yݲ*�ʹ�P��{y#nU��ctܣx�=�L\Ke��d�	і�i�mD�\kKJˋv��N{<�u�gEr�g�(Wx�N���(D�$L�*�b�Q�Wj� 
���c�'c2�Yѝ�y���;:�:ν�:��� �]nL�u�W �3vl����`�lV�0iצWi7:Z�cc����\���A[Z�u���JGu�kQ�����;��C�'��8L�����.[<���LƎ]�j�`u�Ь�]�yv��	�9u�܌I0y���͎�u�yN�=�1Ŭ�����ʵ*�@n�*��N��2y��qP!+U*΋h�&�ćQ��gX��`%�)V�fl�N���T���+Oh�V�mT�U^U�X��
RZ�YU����S�ʂ7s(g]�zb���ι�����Ch�ೲ㬎%ئ�uڜ�[2K�(��*���iT]���l��.��A��6�uEs�����6k,*z�L�/e���b��un�Y�%j����Xjs@nl�\\��BK:�7
j��{V��t���^�9:Ժ����A�z������?G]�����ww6��i&�`  ^��˚b�nKԯ���xG�6��d�Ig�[^t���j)�v�M�A�X0V�����c��;��;�q�;�q�Rَ��q j\��-�h�tŋv�:\���L[T����u���X��e['liS�;I��l�N��pfا��v�8��7_������6s[���mq��v����ӷ-�Bt�aar��P�7iڤ��%;��P��s���-%�֒���p6�f{�S��j��K`f}��`[�8.�ZI����R�8���T-�n���w�˸��E �S.��#��T�a����83"��wQ@�i>�}�`{ޞH�4�"�=��Ƞ�� �+-�w������mm�^P�������:읻8m)c�=��X��g�hxUr�ᴓ��6�&9�'w�3˼�ŵ�1��Im�3"�]��RF�%H!Ű;�f��'������+f<���sl;W���ƻ�b�Ӓ�*���Ǟ��n�(r���;�f���n#�EU)����3"�w�#|�ska�W�}l��+�f�ڶ�Zt��$��(�%�߸�<��9w��&���p�L�w!y{�⬑���ku�ܶ���vLy~�u�B�(�H�� ��mlw�˸��E �S.��#��T*(��ʨ.�o���mo͞�E�T�SR��H�������w�P���RB�.i%(DH�`*��0��b�R�=;��~p��}��]�y�~pmUMS�u�4��*(9���s*�-~�_�� ̬6:��J�[�����ʀr�)䙤�&ir��4�h�,K�����a�ssK[�e�g>��
p�m�U��]82�t�"j�e���{��3K���Kı/�}���S"X�&{�ND�,K�>��:��,K�=���uı,O=������3f]6�q:�bX��}�S�,K���xjr%�bX����N�X6%�|����K��:�y�Wr�ܹ���N�X�%�߿p��Kı;��z8�D��T!�2%���59ı,O>���"X�%�כ���̷L���K���%�by翝N�X�%�|����Kı;����bX���x>'߮����V�*��F�4��3��)�⎤ޗ"X�%�|�}���bX�~��SΪdK��~�Ȗ%�b^����uı,O�&�~�rFɛ�Ba�'��Ѹܛno�m�n6�\vcE[.z�U/���Kı<����bX��:�ޤ��%�bR%��>�'Q,Kľ}�jr%�bX���l35��u���X�%�߿p��Kı/}���:�bX�%��S�,K�;�����*S"X�����eʹ�wf�p�uı,K�~o���b_>�59��@�DȞ}�ND�,K�8jr%�bX�a��웷7n�i�����%�b_?>�ND�,K�}�Ȗ%�bu��5:�D�?&D�9���:�bX�'����	�i��.�3��Kı<����bX�����S��%�b_<��x�D�,K���jr%�bX��}���ۙ�J��,[@  ݭRN�q�k�0��Z�[�[�1�#+�����lG�i�v^�&��$�\���zlne2ݰ�^]a]�T�����\m����vap/m��n�X�v8ٲZ��Y���y�}��dv�nx]�+V�q�ģ���.��g�!r�u��`�١z�'�G=����{����?u��f�c[r]�>�a�O�smU��#x.�͊1Yu-��n��}ı,O�����Kı/}���:�bX�%���jr%�bX���ND�,K�7�n]�t���eӉ�Kı/�{��:�bX�%��S�,K���xjr%�bX�w�ND���D�=��=>.��7&�sw��Kı/ߟ��Ȗ%�bw�59��DȞ���S�,Kľy���:�bX�'���Lɛ!�s6��q:�bX�'�}�S�,K��xjr%�bX����x�D�,K��٩Ȗ%�r��y��3Y��K&i��%�bX���ND�/�2&y�=�'Q,KĽ�����%�bX�}�ND�,K���]��� ��*T�$m�T�)��lXqn�׃��iB(����� �`�,v�{�;�ou�b_}��x�D�,K��٩Ȗ%�bw�4D�,29�>���Kı:óω�sv��乻��%�bX�Ͼ�NC�>�������O"X���ND�,K�<�Ȗ%�d�{����uı,O=��?ni36e�ng�6%�by��59ı,O;���"X6%�{�Ϸ��Kı/�}���bX6']�=��]��v���N�X�%�߿p��Kı;�|��:�bX�%��S�,K���xjr%�bX�y�>����K�k.�N�X�%�������%�bX-��S�,K���9�'"X�%��r�ND�,K��_�㥱�lrs����㗷H�>l���mՋo��S)������-��w�{��7��/�{���bX�'^y�S�,K��jr%�bX�y�=�N�X�%���>ɗ6Cr����Q,K���xjr*��bX�w�ND�,K�<糉�ı/�}����Aʙ��Ϲ���f�r�iwN'Q,K����:��bX�'�y�g��1���H����@ vr�s�����b}�2'���Ȗ%�by��}-�63sL%Ӊ�K�TlO���'Q,Kľ��jr%�bX�y�ND�,lN����"X�%��aߓ���ݻ��.f�:�bX�%��S�,K���xjr%�bX�y�ND�,Jiz�9�.L�f�4���!��5�n����d�Q�q�l,�ҵ:�y`�{���o���M�3r˦��'q,K���jr%�bX�y�ND�,K��=��Kı/�}���bX�'��=��Ss6�3-�8=D�,K�>��D"�	"{��r	 �߾�E$Nw�&���>��,N����3r]�vmeӉ�Kı?>��:�uĤK��٩Ȗ%�bw�59ı,O;���"X�%���g����l7!r��:�bY�Eș���jr%�bX����Ȗ%�by��ND�,ة�b3��DϾ���%�bX�����e�!�n��g��%�bw�59ı,O;���"X�%���s���%�bX�߾�ND�,K��z���~�L���XM<�������c���N�=]؊�"ߎ�{���.��K�q;�bX�'��p��Kı=��{o��%�b_>�O��L�b~eO~��S�lK�����a.	��K���%�b~{�>�N�X�%�}����Kı:�Æ�"X�%��p��ı:ÿ'���ݺnn˻8�D�,K���59ı,�<�Ȗ%�by��ɩȖ%�bw߶cޗ&-3I�]���	QP�u\N�X�%���q��Kı<����b_(�O<��^'Q,EE�/�}���bX�'}�=��]��v�e����%�b{��59ı,N��}�N�X�%�}����Kı:����bX�'����}�ۻ�i�6�Ͷ� <����1�Yõ�pBR�+*�rL�ʓ�5\wH�=��Z#���{x���h,\�-��nn�V�mӉ���2�ڹ�n�xco��?pp����e���4vU�퐈�u�ù�C<@-�9�@B��lT* .��õӵP�.��Ж������[\M#�SȞ���X�iۍ���m����)nx�oz�u�5ps:��k��ػ���d�,K����N�X�%�}����Kı:���b^�dO3�{8�L�f�4�ј����J!#ޗ�,K��٩Ȗ%�`��59ı,O;����%�bw����u�2�D�???�˺ܷww3��Kı<���Ȗ%�by߼59��D�&AȞy��^'Q,KĿ~~f�"X�%��~s�p�5��t����%�b{��ND�,K���o��%�b_~�59ı,N����"X�%��y�ω��l&�K���%�by����uı,?�����D�,K���Ȗ%�by��ND�,K�͞?4�Ihne�Ҏ으��)k�{g].��&|�S�/�\Z�E7�G��%�b_~�59ı,N����"X�%��p��Kı;�~��8i3I�LZ������9D�Sz\"X�'}�G����D���U���K>�;�N�X�%������uİlK��f�"~�@ʙ���=O��Uj���.L�f�4��mD�Kı;�}��:�bX�%�~}u9ı,N����"X�%�מp�f칒�ЗN'Q,K �<�~��:�bX�%��S�,K���}��uİ?	�>��S�,K��ͦ/'#�A!#r=�p�f�4����T�Ȗ%�bu�59ı,O;���"X�%��{����Kı=��߾\�Ks�����t�7vu�����v5s٫��#{���8^wH]�ww3��Kı{����bX�'���S�,K������%�bX�߾�ND�,K���e�a��̺\Ӊ�Kı=����X�%��{ﻜN�X�%�}����Kı;�����bX�y���]6sp�N'Q,K�������ʙ"X�߹���c���������wM� �m$�K	�c�6�[��O+��:A`]�"���s u�Ѳ�}!O�!t���W��{�B!d��0bXBD���;%��*���AȐ����RwP���QlW0� �/0 hrd5�Ra�x�t��#אT(C�w�t%�/J&+��� z��|�^���T����?bwϽ�Ȗ%�b~w��S�,K�����2��ni3v�:�bX�%�����Kı:����bX�'���S�,K,N�߽�N�\��2'��߲Kѹ�2�3��JD�,N����"X�%��~���Kı;��{8�D�,K���jr%�b���Z�p���FZ��� 1
���\�Nָ{���.�!R�]'��e��V�����q�ı>��"X�%��~����%�bX��ϳC�H�Q2%�bw��59�L��<�o�?3&�B��8�D�,K�?9���ı,K��f�"X�%�׾���K��<����،�f��X�#d�G*���&h�/�}���bX�'^��S�,K��jr%�bX���=�N�X�%���N}2��!v����'Q,K?RD���S�,K��ϸjr%�bX������uİ?G�������_���Kı;�M��Y��ۗL�8�D�,K�>�Ȗ%�bw߼�q:�bX�%��S�,K���xjr)�L�f�m�n7UUCN�j�\�ݽVDǮ�Հ�q\��g�RZ����g�w���K�2&D������%�bX�߾�ND�,K�|�Ȗ%�by��59ı,N����.�f曹���Kı/�}�<�bX6'^��S�,K��jr%�bX���{x�D�,K�Ͼ$�!�����q:�bX�'{�S�,K��xjr%ڙ"w����uı,K���"X�%�מY�R����2��Ӊ�Kı=����bX�'���'Q,Kľ��jr%�bX���ND�,K�&��fI�d��3N'Q,K�������%�bX~�Ͽ?3S���2&D��xjr%�bX�w��S�,K����|`v�h&$H:�w�������d�m� m��;u�j%�X�.��6,�l�;պ�4suòƱ��g
��mɰ�����n�1��9�Ɠ���Tu�C۵�p<��t��-]����b����\�Wf�x���z�+R1<��X�,vH�]�!q�ۀ�[����[�뜻9�b9�vm�K��o�����:-�Fɰ��Emɸx���q���Wt�VAns>83��2�mͽ'�Kı/�ϳS�,K���8jr%�bX�w��S�,Kĺ��[���&i3K��~)ӑ������%�bX�{�ND�,K�=��6%�by�y�q:�bXL���٩Ȗ%�b{���a�͹w&i��%�bX���ND�,K���s��K �,K��f�s��ı=�8jr%�bX=�|m�sk.��f�N�X�%��}��8�D�,K���jr%�bX���ND�,K���Ȗ)�L����*�u"�$��p�f�ľ��jr%�bX�{�59ı,O;���"X�%��}���%�f�4�xx�`����'��M��蕦��k�]]9�Ʌ���h�K!v�~=ߝ�7��,N����"X�%��~���Kı<Ͻ�8N�dK��>���Kı;��9�vf��r����%"X�'�}�S����@5{P�� N�u��>����%�bX���S�,K���8]NDȖ%��|���7�4&k��%�bX�����N�X�%��}���K�gu6'��ND�,K�?8jr%�bX?����.��nm6��q:�bX%���}u9ı,O|����Kı;���"X�%��}���%�bX���Ϧ\���dۻ���Kı>����bX�j!�~�juı,O3�=�'Q,K��>��r%�bX������;*L�#{��'d��#fN�y��4�W=3����Y��۔�&i��%�bX�y�ND�,K���s��Kı>Ͼ���΢dK���xjr%�bX����Y�����3N'Q,K��=��8�C��DȖ'�~~]ND�,K��Ȗ%�bw��ND�DȖ&"wO��U���I��4,гB������%�bX���ND�� ?�T1�D�&}���q:�bX�'�?^����ı=}��ѹ���&��uı,O����"X�%��~���Kı<�>�8�D�,K���Ȗ%�D�;���3ws�st�uı,Kߟf�"X�%��y���%�bX�g�]ND�,K�|�Ȗ%�b~!�������ṳ2cI����!!z˯Y�ڷQ��f�f�m�2���O�����%�b}�~~g��%�b}��u9ı,O}�"X�%�z����ı>�'��sr���sw8�D�,K���ȶ"X���=�N�X�%�{����Kʙ"{���q:�bX����ߊt�C G%=����L�f��{�G�,KĽ��jr%�bX�g�{�N�X�%��{���Kİ}�|���3Bne�3N'Q,K?Q��3�3S�,K��=���uĬK�=��r%�`~�p��-�XHS��#Ҁb"a	�O����I�L�f��/�QF�$	z\4�K��=��8�D�,K���Ȗ�b{�59ı,N����"X��f���7�
G)S��)�B�Jfr������խ�]!�W��$!`ڵ�r@�g����q�ı?3�˩Ȗ%�b{�59ı,N���Ȗ%�by����N�s*dKϡ�����nɻx�D�,K�=���dL�bg~���Kı<��}8�D�,K����NDȖ%��~_z�n˻��f\�8�D�,K�>�Ȗ%�byߜ�q:�c�(G"dO������bR%���p��Lʙ��ɾL��n̗4&i��%�bX���?'��%�b}�}u9ı,O|���"X��2'�~tjr%�bX����~��䰻�rfl�uı,O��߳��Kı>����bX�'���S�,K��9��uı,O۾��w�^��{��qo^���` *��8o���}�^m�a�vK�R�dG)�n��t����5��u|��f��i�=�`��<W���&�M�<��S��Ew6i�W=�f�
�U�j�9Nz��c*��
������ȳL�x`��!�n�w"q�
jH�X0;\��igX����o�w����%v�v���.???q�G��h2v7�mٻ�U���+��35S6e˺B�wr��D�,K����Ȗ%�bw߼59ı,O;��uı,O�Ȗ%�b{���at&�ݙ���%�by��59�r&D�=��}8�D�,K�??.�"X�%�����Kı<�|��l���v䛸q:�bX�'�o�^'Q,KĿ}�jr%�bX���ND�,K��䚜�bX�'Fxy�Wm��fm�uĳ�#��٩�Kı>����bX�'}��S�,K�<�}x�D�,Kϡ��ѹ���7s��K�,O����"X�%��~���Kı<�|��:�bX�%��S�lK��;�}�6���,�<�v�o%ۢRV�!�IP�q�t�6iIē<Լ����%�bX�y>�Ȗ%�by����uı,K��f�"X�%ʞ��F�Q,K��ɾL�2]�.�fi��%�bX����x�B!����؛�����"]��2'���S�,K�����bX�'�y=��7!e��乷��Kı=�}�ND�,K�=�Ȗ%�bw��59ı,O;�N'Q,K���}2�݅�6�7��Kı>��<�bX�'}��S�,K��9��uı,O~����bX�'�o�ˆK.ܻ�4�uı,O|���"X�-��~s���%�bX�}>�"X�%�����K�7��~C��&{j<΀��`0��� �w=�Җ�����g���v���~7���{����>���%�b{����K�,O|����`�'����I�|n��swff�A$O��b}ı<����bX�'}��S�,K���}��u�,Kϡ��ѹ�s.���uı,O}���"X�%��~���K�@@�B��J�D�UZ �E|z|XȞD��Ϻ8�D�,K�y�jr%�bX���z˳7n�.nN�X�%��p��Kı=��z���%�bY��������K�芹����Kı=�o�?&d͙.�fi��%�bX��{�G��%�b_~�f�"X�%��~s&�"X�%��p��Kı;��)U8��Z�QSR��MU"x۵p�q��ci-����s�Y��10������oq��٩Ȗ%�b{�59ı,N������bX�'��ϧ��%�b}��>�r�ܷww3��KĽT�ߺ5:��9��,O����"X�%��s�q:�bX�%�����Kı=�|�\0�Bf��4�uı,O|���"X�%��~s���%�bX�߾�ND�,K�=�Ȗ%�bwޞS�K�m�s0����%�����q:�bX�%��sG�,K���xjr%�`~��=E��}P�Q?[�Rjr%�bX�������)���%ݜN�X�%�|�{���yS"dO|���"X�%��~p��Kľy�>�������ݵ�lw-��0�3kŻv+��iq�:���TN��Q�6�$��q��bd��=?
��V"O��d���Ɠ-�h&�ԥ�>����Y����� �J�YT8P�MA��w0�]�<��y��q@<�]�ԡ�ʎ��6뺀]ڊ��P����jaN��P�$�[3"�_{>n�獀Xf6��$�𻰑I  <��xM�!�g�U^�I�y�~���Q=`W;| >(CҀ���B#��De@�B���bgjRY	 Nièb��HBc�W�Ә�j���tJI�)� #�o��RH���&�F��cUUA�m��    $ ��"F� [��� m               ��m&S��=�؍��l�l���[.��ڮq �5��cTٶ�g����@b^����V�;Rh� f��ݤ��gu���f���\J��U*��K���k��)E[j�s�c��6����IZ�4��P㔉N��p���`x�Vq5+���R�O..�ck6�6`�^#E��a��SM�,{�@nҺ�#;������1��ѵ�"�)#?t�
} mɹVe�V��Bt-��7[ulk[���'
������$��N�5 ۖ%�Zn�#tdk�-���q�����y��3��ʭ�B�b��w6�`V�(�ʵl�����+�W֌-��2��ghxy�g�iU����m�{�y�� ��zݲY�r@ "m*�vդ����0&{�[�]Nݞ���;uv��l�U�;Qc�Q��m��eAuaI�3�ŧ���8g6qm�5kW/@m�W&�Z�4gn�:�X봶x8uZ��q6x�l:n���%1˵QnY媃�����o-�n�������m�R�y'm�ut�϶e��UX)V�fl�;��ڹ`T6�q ��yZ���U�3�]�[M�bYR-�� i�$0�I���d�t�s)��.X[���+<�f�{g�m�6�p^Hv��G�������8	� *fMT.��������Y�v�Y�9�����}:��s�sէi�w�ڌIu�#S�nm��;<�ij��KH�DҬd&���(q�b�Մ�s����2h-�un̝]C.����������M$@G�?G�P��g���z��x.��)���~w��|�������wX�� �=ORT`���,.x'���7W`ݢ��o���1��}����a���s�[�Ml7n6�8%V��z@�mo9��h���6mD�����#�H<��ֳ���gF٬��rg��糹g mv�r*p��W7Y(�#nܚA��F������Z]%�.l��vi�Iꈷ�����S;%�k��B�whe8�T�D(�K��F��w�M�Tɦ���g���Y��u �����o���r�$\3�	'dL�$a�w1��_PH��m*j7R&� �ި��i-ii���]��=ՙ��'U
q�`f^ml��w�f�2�}��)I�N�J\�q�%w{À����̊�c��2P'MPƁ���������nz3���=�]���s:81D�,��.�m��~������]�P�c�v�R�'*4�3�J����?::���@ �����gk���|o����g��<S�"��U����5 �*�{��`�*˻�n�9��$�)lv��w��l/*wq@;�]xFUE)���� �ʀ]�P�y-%�j�h�N���P.����u�^�st��L>֦�qy���JT�nH�� �z�ý� |�=���X]���|���U"*�N"Ul�K���j��K$����I�jd��
���)It�T�� �W���f����UT����;�Œ{�}-����:
������s*�ՐA��vv��P��GT� �e@?i%�+����׈���`_�&�5��	 ��%�,K�i�n�������*箋�lul��t��Ul���U����^e@9w{#����DU(���{I&�]ņ�3ި���]��U�U"��˹��/0�{V@;������GMF�u�������ި�a��_r�]��p �Ub@ `������{	?`���M��*�;K`_kyV@7ܽ���y��7}0�ۣe�����5��68�V鬍':Goq-�&�쎢��G*R�9J�Tp��a8�����y��ݰ���?d�Lp�ST7��fmo���a��@;���]x�y�Yhu(L�9%E��ɰ;��Ii7�V@9�ͭ���`U!B��*�{X@'y,�����/2����U:sCqER�X@7w{[ �ʀ;ن�~�� 	�=�s��ݷ���u��  Nk�GS�˓^�Y\D�*��et�\��H���N���xࠡgv�um�Q��v�����ĺ�<U��nQ��n�nD苶��6;m��B|���Ѫ�v����aD�� 8�ö�Z!�dj�<�Q�s����-��$5�rc�j󆍅b�]��ٿ�����{w���p;�����w)�=/m���pq��V��W+�{S����GU!p���o[ �ʀo�ekIF�a���U�`H�ܑJ����@7ʲ�W�󷵰9�ie�����@���������o;{[ �e@7�ٹR)QƩ�G�ˬ ����;�P=����ǰ/)�Д:u4�ۼ��Zw�V��������e�붰ձ�iǝ�y�wl����%�B��V5����olJ%T�$�����Ր��@7̽��3	�U��NT��`r�	�\ZI-$�������6��eO��Zl�����9�����ܯ��k`y�8�V@:��X��R:�$n���ݶc���;p:�ل���	5�'*-����l�rx����z���~opQ�pQ�Rt�[:�v�
�HK�q=ve�XB%nt��QJ��$IQ�]a �*Ȁ�2���y���7*E*8�:��9�� �.��;Ơ�Y �i��P8���T6;���Oo�ݟ�����bw�g�"�V�*W9_���
�T�p�-��p���o��|����f�t�!B��)�]a �*�����1�' ���`�aLC���r��zf�<�a��.�L`^6#��9�9�!q�t�[�;X@7˽Ѱ1�?m�{X@-���UQH�I)�lwٵ�1�8�V@9��ğXH�#rD�E�1�8�W��v�@9�f���,�ۨ�����pu�|� �^���崵BY�!)�IT(�>۲O:�켧
��T�TN�U��]�lw��Ր�i%�cm7��PN�J��*�θ�2�2!�-�'�-{F���sf��4#{fN����<�o�X�;]'1ݽ���OQ�	"��}*��X@7ܽ����6S�)�J������o�{[�v��dt�I�"����k�w��1�8Z��� )�I0ٴ�Wl������r�-�I�j��X@6�]֓�4�@�B�����Ds��m�  ,W�,�WM��R����;��֫���y��-�j������,�ō����z�����J�΀�z����W�7g!��u�Ss��	�O+���Ȼ�P�q�kI��.B��[;�ƺ.pmD��;x�;]�YLԯjv��{5��X�c8��7�7d��7OA�TP�?wg}v�ۨ�Kc[��.��:±����/�k�$Vť�'N�)H��DnH�����p���o���e�l�fl��4�"2���1�7ʲ�e��ŭ6v�)�*�����Ƞ�������V@;ҲӔʎ�MF������}� 4��{P<��*�S�!	"�}� �j��wk`s�{[k�Y��ʟ��"�N����DLrpm�ݻ7�Z����(;h�r$�M'�m���u��Ƞ�b�[�\�]�:o�9DUU/6��~i���+��F@	��\�;T �û=��N��d�b��vy������
�I��I3}�$����o�d9q@8�qG��H�Ql�ߝ�r��ؠ�k`e�3nR��U#��¢a|�Pw/k`,}� ;�w"��$D�l��������s��th������f�ٛ3�5�n�m�~W@7˽������Z �<�R�p���8�;��6;� ��f>˸�w�l*�S�!	"���o�d;�nu�x�dr �1a��i�!�� 3�{� ��w�9�S� Fp��_� z�D�or3(�Yʀ��9|=	$��"�H1HA���		�ǭ�P�H�x�07N8�F!�,l���	 ��v�1L\h�z�I�%�Á$
$F�X����F@!U���,�F�Oz����끂��k*�(��E� I��$"hE��$=m�q�'B�^��21�BO}�0`H�	� �	���Hz�E�p=�! �9zȑ1� &�h�`v���}����u�"��(r{��T )��?�]" ��@#��'������hV��M+m:{��}���j(����wn�ꖣ)�BUF�T6]� ��c��V@��w ��)�U	A÷ �v�p�GG�����Tn����#sv[��{�w3k`˨�V@2���e���7R"T�`���U��e����ߖ��M��{�n���T��ܯ���k`2�|핺*$j���2�o�{[�����h;ʠH���FH� �"B
�! �#��,��"$�0`�b��,H*d�"��I  � �$(T(z���w�W��I4�I�6���~ͭ�ay� ���� ޙ�wt�ql�yw<]t��'<m���*�g������٢�GDa*U=�-�w.��Y ��P:��6����S�(Ԣ9)�v���I�2�sכ[�gY�S�-$�8���T�*������(ﷺ6I��c�p�;������m�
��.0{X�n�B��5���x;d���t�03��v᭝�sr0>
��� ��Οk��z�Y�h  '�H�y�#���vn��I�&F͜�X�6[���7��-^�/'M��'$����X�1q�
q��Cu��O�;v��b�����1���`l�C�n��E���+�i��[C̾1fK ��WkGV�i�n�ݮ����09u���1��������0ٻ��w���tv?�{`8�W_��� nW}\d�]�+���U�5�ۈr7&���*|���i�|��203a�s2+j�ݧn¶ػf�sX���gv1��5��ح��)'I�\٬��9ۆ�vN	��v�wE�ݶ̌s�l�c����G}4�j�,�n�\/Ƥ�c�����br�S��My�ۣ�%��@����-��Eۘ�F��Q����a&kw5�L��gv1��A��@Ra���v�p��=��'�Q_��Q�@�/Ƨ$c��g��J.�6�{��kt<k�ry�XD�L������br<���S�1͊�v1ܗ6�M�
�l��u�H���c��'��d3e�1���Gn8"�v�r%����\a7�#��L�����}׾����{p�v�c6�ƅ���l�w]��;ۆ��1ͼ�YݸV�j�!�n�C��zjrG�5@	U���v�
� 0P�o��k��bf(.л`&�	3[��91C]��9ۆ�����j�6�K��5�����w/M{�1��p�v�b}�y�Q6��n͞ 9]�n�����1[�}@�ev�%�`s��n�dc����MZ��.Շe��r�ԙ��`gsX�KQ�&��i;`�ɬrdu����1���8{~���-+`��;饁2k���@N�*���_�|�N��* SN�[����s�gsX��a}~X�����	@�%H5P��Os: 5:�Ȯ�ۉ�y�nͻ�
մC*�i�d���c�����3�h+`&�	24���&Fɬs�����<�I���m]����2k��r��<�A��ݔ��l;L	�X�n������5�틲�%��r��w#܌	�S� m
����ӻ�����-��,[@�
��n%��Sγ�nC�k��g٫��K��'�����p6�\����ys���R��V�ԪE؞�vƶا/]jnD�w�#E�����9=�N�l�F�U�a��vsƫ��k�įN6�t*u�X���
g=��]��2�H&vXL �,&�Vڡ@W��(�Y�ζd̲fId,ɛ�hd��uV��ɮ�n���p��s^��G3�a���??��L�	��v�p��"�,���S���`L��;p�w5��o
�ݦ��-��&Mc��k���;��ݚu���D2�����5���;���5�1K�A&h��5�5�vFdׇ�p��
��#/���M�v����{v���\XOb�9��JJ�UTR7"�np;~�K���Ö��k��1���ݖ��-03'����h�j���Q���D +(�!I�@�um�<翚s��4<'�'l]�um�;/Mgr?����6o�Γ��l��i�ͦ��[61����5��Q]w���-"]�SS�ɺ��5��ٮ�3���AԐ�T9T>w��=�����Xy�-��:�xس=��f�U�������e驓�lt;��Z����a��&^�}��3cd�$�`��E��������5�0_`�'��b)�-�����O��|L7m�����f��f����Y��Fh,�ݒ��m�&M|=n�w�ȷܸ���o ��ࢦ��D��g*�:ZkՃ(��Q+tX�v���WV���zjd�9�52k�ܼR�,�����횝��2Fɬgn�	��mY�lYO��u�2kۆ���wo
�۰-0�n�EU
��|�;/ƦO���w@RZē�I+��{���
�*mn�i���l`L���BE�%Y$��=s��v x�yݼ��7l�i�
��&K\<�sf�)�D����F2o���\̈�$�n�I]��������������|�џ�n�)�[f�Ml�lCO��s�jL�6�b�E��o�����c��L��;qK,��v�횙5����+'�����oW�����䐄��2e���������U?��%E�9���:�:?�mxfC!��c��J)�����"#U!$�'�� H#��  ��G @�B �g�j�bA��R@@# ��rU6,RA�$b(���(H
�� *8Z������ ���  ���(H��"�F  �"� `
*H��B �� C
�.A, EIh�&P�A��Eꋫ�����a�����A�>�������o�|A?�Q�~b���A2*;���p����S�DO�����������(3_�E�7���Z�:������d9�
<4���3Ҽ�*�9׀  ��������?��I��?����?� A�����?���O�����g���!��!����C���� ���?̈��T������#���P����O��Ȳ���t����������9�۽A�~����T�n����ӯ��M�D(�� E�����!	!"I$ ���H����H� A?��� � H��"�H22!",���! "�",�Ȳ�I6� ��B H���  '��"Ȫ� 	 $��"B$!"H��,""H* � �",��*�
�2)F 2* ��"���(� ��
�B(� +,�) � �!!""#"�(�"� �!"�
0���H� �2����(��`(�(�������`�E�T��@ (�P ����� ����"�V(�
,U���� �"�A��D��(����`�`���F�`(�A��Ā�@
�R(�*�D (��"�
� �@(� 
������ 
D �@��AX�,P �D",Q"(0 $X�Fy���Ɠ��)�<���ƽ���C�g����""���;�����y�?���������R��?c���?�?�i���t'�����! A?���MO����_����	��7�w��N#���o�9�����S���O���~?���;� � ���
(@�-���_ɓ�����?��ާ��#��K ��G�O�" �?���Τ?����	����_���SÄ��C���D@A?u���I*~��G? �#R���PwB��Blm�A��8�����#��Ґ��vt�?���`� � ����b������?��������	�����Al��������/��������� �?�	�����P #��P�<?�����������/��_�C�/���	���R��ie���&��%��"F��O�S��ӏǰ@G��t�H~��� _���W����O��O"�'�úhp��������G� �@G���q���޾A� ���s��v(�#�B���^o���9�4?��ߊi/�|���rE8P��`g