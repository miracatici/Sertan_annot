BZh91AY&SYX"���_�pp��b� ����ak� (���P ��) U��QP������� 
)*�JI*�)J���@��R �$A@ �B�  (
H�� �@( �� @ 	(��( $Q�   ,
@ �P�(b }��b;�S��0q� {ޔ���K�@�1 � (�}5�	5� R�ZUfk�T� �CJ���R��
&�j���U14�CJ�m� Ӊ���    }� @  
�(��� �}5�����yiO\��n ������1w4�dWs�]�0��@u*��cc��o0����8 ���!�2轻�����=}��\�}z_|��˞Ξ[�e\ ���    �(e� �=���{�{3�Ҿ۞��� ���˺ڷ9�lq�u�̣ �9o{r^{ z�`���� ����t�{����7��� ���a����\Z�NAǀ�|    �I@Q�� }�I��7<�绔90=���
��@����X>V{p7z ���0�8����Eɡy�>�:w�J����<��q�ڗ6��y���L�Kv;�s�]/y��xT� @	 (Š ����냌|�\�t����Tn >���7��{ŗ6����x�����*�wV�c�  ��v�v��(� ,�����G��:b��7��{�ϱ�9>��<�K�@       O�&��U*��4�   �ODCRT� @ ��OǪ�J��      D�*��d�F  #  0EO�&�m��U�@� A�� �!T�4*{Dѩ�4�Fjj�ȟ���?������퇷��:��u��QU}_� 
��AUO芢��p
�����**���EU�����"����?���������_�o��۫9�J�����ba	BP��P�M$x��	BR�a��m��C��&�H�0���#@d8	�a��jC2QD����N����05u��<�0r`���a97��k����Z;2��%��9٠�jv���S)]	��$j���]�Uw^�y&&N/3�(MBw.�؆C���E:��՘xAb��s��vk{��/BN��j8��P�7�B��T�h�E�.�2p��8c��]l��3h6mٜ�ё&�;��g�Ӥԇ(cElk	��%)I�U�ĴRZ�;ɞ�\�G��s1;�FP�ł�:R�x��)�=q{}�­Z6���ۼ�#�Y�v���+9j�<�ʿL���Vګ�u"M���ѫ ��1�'#N6�f�4F4��8��b�6i��r*(�bCHMAʢ:��	!�!������0�V��`�H�j���Er�ğ3���.Z��� ��2C;�@��C20�\��0"ˮn���t:\���9h�u�^6/r�m���]m�)̒8��X��
��m�;��I��SLL5=�发YJ	&��p����J�JPs&F=�22�6�͜-�J4a��� v'#a�i��*4dky��������Ĵ���ӽ܍��'3C���>:�4e�l�ﾇp��b��]o�u��'������s���vqv���N�N���s��w;�Y;ξLZ�	`�>�W�![�룮��w�q�9�Ҹ���ɺ�ꜘ��O#x�C��ȉ7w�WV�Q�1����A�����`�%L73�j��306���:��;�&��÷W�2&��<9��`t��p�9bn{�&��v'D��s � ��ɦ$*V�+),�"��m��F����}�z���$��S�N���i	�I2Sm��!��Z�B�Rb)�x�[�|�g$���h|�$W`�)10�z5V�X�MF���-�rR����䆼�����ӳ�ב�;�!(rwY	BP�%	����,��dt���:<=��k9��2�8F�*�8��kq�[��d�d��&����:�e1d�K�"~bYײsYb�	��`]Bw	�'R&Bw���՚n�����?:h�˂&OB����]���	��N]s��ƪ%�$�
�jP�&BP��yt�y�;�'���N�[Ow�A���V�.FнB��(��H�^��C����/uh����<��JFX�`�5�NBd���GI�p��a���Qu���U��W!�z��:[�Eԅ������Ӣ���NbBwe4�jLL�H���f���2Xv�qy�rd%'d�A�^`kw}����0�u.9	Ho �4owy]�7�Y���4�	A��3ս=��'Qo\���C�Q�v����Y���Rx�Z�u�CYc���C[h���o�F�79���@hE.H�V�R�J��Χ,^����:�L�&L5ks��tXaĜ'F�sFНBf�6��;��I���q��n	�H��J!!E��[V���;���P���i7��%�bu)K�t�*�{�W�N�D�$�#�o.�|����o��;zN��ut�������	H�J�5q�?w"9��yǋ���x1Z�.�E IO��P���.�:6��ظ�fb�z��hS����y8�fq	�.�E�$�P&����N0gDRwf݆�\�����^������S��5G(;�<Ԙ���x'!%�qtÖ�NN��5�.BPf�����npĝ@�BPOdR�٫F���³BP���u���q]��f�N�Ih�!"��1۬����X����uu�{ѷP`��]�'%�#Aǽ���1��F�����V�Ru�:\�e�a�ӑ���8w���L�&w7wX��(6�CYd��|��E�H��c�j2�*xfsi`��K�0��!"��(����F*u	�c��,s�#� �3.��{՝/�Z�T&��u	�L�'[qz�����:*��5t�CУgoG��,tfdbtnC��H����g'���|M����rd���s2u�n�N�����˱(JItK��M�	F���S�Z�$��>�3�X�9���T�R�%�i�(N�(Mfi&,��(MK��Ų�0((����3b�DD�5NRv�2��D��Ƚ��)�(F�P�v��L�99h7��{5��F2`�&%h�T��=DQ�Iq���YO˙����QN��%	By�%'!)�� �0��BQ-I���(v	X:u�k!:��%	m��m�t���f��w7���_���8Ì�h3f��h�7�dR	J҂�HN�A�M
��~�g���"��+H���kQ3/���h]��,�Zs�ư�$I�u%#�f�9����gIզpXp��.BS�I���l���^w�{و�5�����c���4�7�����-e���%	�`�hv'����Yb��dU;�6:H����� :�3T:��㓁9b��0�SW�)�����ђ�A$�k�j���(J�N�̪����V���V�S<�k#LMڟ�������G`d%`�ԛ�������[����F3X����x:�cXj0c!�2qr���lj���S�D8R�Y�g�4f��Gv���J0 ���%óY�2��6�.9h�ѷ��������7�&�4���{8��a⩧�����K����pY��e5Bk�i(1&��BVqx�)y>ԦZo8�EA)N�Q4��/����	OnP]�An��-`hr�1�l1uZ�ߗ�����U���+X�������Ԅ���6٣|��}	��+�8U:�k;��Dƭe�����l9bHfB{�������e:bi&W�om��h�M-v�ʳg�7'!,to�NXi2q5γ�_2�W�:�8վ5�I�K)ASI�V�@wR`S�٩q�Hy��@]V9��QCE,��-'hN��CPNJ�%�b@�����ї��ZC@4�@��"���(������	�㓁>kbP��w���6�]o\�Lt���"���iݩ���ʧ�K�GP�ړ���jj(���6U�(��(1�`Q��双5ִrZ���;���q�|ER3�F�in���r5Bt*�D��0��R�P%!��rl�-�����5�Q���Uݫ������/M�ъv�y�Ve�;�����R�����J۸Os��2���|���7a��z�Qq_0��WQ��-X�kcJr�	4����Ms.��H�����9�]��.Z=/c[d�v'��`c:uP�� ĺ��{�t��0jpl�g���o���'M�����^�֠9���<�����2���3�0J5��y:�I��&A�d�k02c�2����[
�X^;k#��h���cGrcXڃ���Խ:� 0ܸ���ĕ�k��\��!g��_ �4'���p꬗\���m�	:�{<�W�<:|��������v!���}\�b`]I���6�Z��@QQ}p/
uek�I����:J7KPd'��K��%!�&&BP��rC31cq�r#�:ܹ]��-����h����"Z痺�\��.��媲��pJ%H"ʇ�pd����3�^V�P�\�<D�LIѣ.�ueW��p���.Ύ&�)|r\s�R��ē)���Xz�-�Y
��(>&�����y�0x����(IԑԘ����Hw�	NY	p�4fEW���t߮�O����Rʜ��S��aPL]iH�T�wU�r�
�&]bMz���r�6n�D���&u.���u�������N����]9t�4�i4%
i���W��S3�\s������3�%� �L5��A�q�&��Nf	�v:T)ʔ�A�M�t�bqB�u���WI��)z��e�q�JˆB{['ZN��4S��Bxf	C�e��A��J�(JbE2V�,�/8�(�̤�P�T�P�D��F^ALQ�����RTjU��ݝl�C2LN�0�qr0����U5%�Z���K)��[h��IpM�6� c>N�,��[ӵ��A�	R��l��K�T
���R㐚��P���z���:�$3�Oa(Ou�r��lC�D�F�2tY`A���`����dh�W��F�4;���=��`�3���w	A�*��8NBP�'Y�Z6��ݺ���`�u:��%	hƁbn��R���块o
M�����D�aw�w٣w�۪��8;\�����̓,��C2ͥ��Q"A�ɅНيv,��%*;h2�`Y	X�7�&���ЗYlãs���ij�C�΂]�EW*"�(�Ȯ
]�P�2M��:�'K��r^���!2���bL\ۺzSci���SSI#>f!$�&��#2r�"d���N��23�3;�N:��o�IOA�V$���N��*^n x�W�g�׿���:x���  �   3�Hm�   3�@hd
P`�`   9�  R�  ��   H  �-�6��!�@� p���A   ��M�mp����h.�ܠ]����b%�J�t��vevv5�mv$N�I�I# �o@[�u*�6�8����i�#��kj�  [u@*��7��]���VV�J�l08�aZ�R@j���tJ�*��O9zD�@B�UmT�|pZ����*�'�:aF4�	;�;��m��.3F*�%�[U�p�g@�6�j�[m�Op[�������[��4"q�H&�H���846��JV��++�u@uu�� 僂�UWX .Wm�����&�b�I:�]~����흞�Rl���5Ҫ��p�N�\�;eV�x�yn�K#�䶮�\ڬ��:�2p����m�ew-gA�Q\h�dSu�����&r5�m�H��[%��rm%�����(UUL=�8 �M��:���n�����P�����6�E�qm v�i6�V��O�g [D�s�J�  8�n�m��Z�m��\I�]��%    �u�o�]n-6��(�p ��}m�3glձm   m{ 8m�e�Jj�
�9P,HClg�Ai��eZ��s�j�f����p��%�K�Z� �!C#�MqM[   �\��Mm�?T��헭�� �`� �kkFݴ��#��#�]�ئ�ٺ��۰�U��P��E�=�55X����dHs[HM��h$  �o�   ��H�n�,K��h	�m���:�)'-�8����m�	 �b�-�K�ݶ�  n��� $  a��ŷ�hp [|&���n�h-���˷d�j����*U�v!����1Su VR�ͳ�$#]]c�T�=��	  �`7m��p-��\��  ��,�ު�U�nͮ��s ����W��H�x�5Tkj��av��n�\m[6�	��[K��	����`�+����m�6�I'��o0ր d�f6��f�v� o�{Io{�$ 6�*ʵ�R�u���#m1� ��[I����!m�	$$�����d�� ���� �[@ �u�      m�kp�� !!�v�fݰmm�m�ŷ���H6�m-��pj� ��   6� r�n�ph8 �  m�p�8 �@�a�� ����A�� �  .�j��Ҁ�U�W�{��`�H q'm&�@��h  ڶ  8��M��*Ҫn�P��j��6@KU��P� ��M�}�Im��l҇,4�l-��@���� ��06�m�3l�m-i7[@��3$����[��y��݆�4�c;,Z�Jp��g6��+�����m$t�fqU�9�)I�����tS��hsm��KWl6�fε�l�` հZ����	��	f���� ��Hm�[@�m���j2ͪB�mʭmW[l�
�r�H� ��MڂA�)�Ͷp���� ���NkZ�(L͖�8�   �Im5�[RH��E���l &̣�<�p q����� �`� 7m���[m�m�-��� p  7m���   ��޴ȡ#v�n�@:j�8� m�kX��� m�Z��Ͱ$    6ͱ!�ַ�I��hp 5� m -��I�Y%�� ����k@ ���I���]0��& �t�f��8	me��Ѫ�����U�44I:]�`m����` �����#�d� m� �F�Ѷ��-�m۰8mm�d��݅�1���t���]iQ��4�:�l6��v ��A��[�@l��m�N����	�v���� [@6�8 m�m%�� <ڳll�8�۳��m����5���L�Z�����7�vHӬ4�[��[m�� 8�k��  �m%�mní�n Y� �Am�N��{��w�::U��yYvZ�	V��[�� h���,2ր:G 	Kh���4vN\���UJ�D�Ig6@�jW���]AH��U]�z�R�3����� �֍���F����\Q�$Ud���'(�����UPq�U9n۵��` �^�5�Y�M���6��R���̪��A���$8�V���6�v�ih�ѵU�K�d6a��r�h��Y!�d��[i �8mH` s�i'9�6� 6��m2�z��q��e�m��ګ`F��`,6��!�Mn-�%f��  g�da,�9�����$��{�M='FY�L��m�k�p����]�m�;Wgx�v�-ʪ�6{���<�үSI�� ��-�8�<(��H	@��R��������(��-�ݕt]�*�@U[Sq�%Z��*���@9���RAR�(n�Fu�-.a��������pY�7C�P�ڪ�W��%�k�\@Vբ�   t�k��5�P�m��'@	 m��mK��:M��`�� �e����H �ߏp���o` 6�[lp��h�  H6� m���-h$�l-�lN�5�$�m&��#����]m"͑��f� pr�UP�(M�
�
�}�m�%���]ml��s�	�&F5�  [E���   6�@m��lӒ$Ӏ���h�)��m�m� �l �a��$�" Xl�'YE#���7�.���
�V��j�r�����   Hm�l-�  �: G�N�7��'Z�Ā� 6��V�m�[@ �v��� �9[I%V�v�k��Č��`   n�$�6� &� �i6�t%��n���� 5�m qR�J���.ԪpPR�(6�Au�,S��WD����Z�6�2��UZ�.� m-��6�-p[F�u�u�9����I���$m&�ƲIIl��/P� Ӷ/E�}��P�^�8p8�m&À���� �/;�X�KCne�Fɰ�b�vXyڥn�wm�UZ�V>��9Nۓ!�%w8*�T�++@U@ Uj�H�x����m� �+ga�׋>��se�`�8iw.��9����ä���;V�8�!q�'ɮ�l�=6��>�·vZ֬�$q� ��<�����W.BƅR����9#�lX@��L�UN�VԦ�8`-� ��ځ9�� �n� [FҮ ���� p6Z�I�����	 Ύ�b�&t�@ �  ��� 8�gi��A��mo��O�4F�fsm�m�@���֤    �b� [Am8H ��8 	�� �v�      �h5�m�6� ��]6��mt ��  �^�m�`m� �M�)<�R�>^j�m��       � A�$$m��K�it��Um�ѯV��h�hIoU�a����&�6� 8�m��om��N�A �,1���� $n� p8  z��ض�m"E�  ږ�@�[p	�   �6�@$  �` � �@l ڴ�  -6 h   ;Z�m�� ۭ`$�l  ��h �u- ���[[vKL��WeTr�UUP��P�/UW����حHR�ֵ� ��e�:�[@  � m����:%RZ�V���U��������$2$��Ra�ڽ0m�m p  e�R����T�]b�H݈ �5�I��,�mV9�ޥ��մ$�W�
^z�UZH��V��`�    	0��-����ۤ�kn�ݖC��m6`Ø�����;:Ѷ���rPֈ*�mUJ�U@WUJ��(p���*h$5��j����5q�8���k/g��]j��̫tF�evv^�V��Z�f�(��6z͹KE�=��m�f��g�e��X
��[N l��k^�D�	l ����� ! ��ԫ+k�m 6� �      <m��h�ɶ���7oxx8m[h�6Ѯ �Ͷ��: �b�@�@��X    �   ��m��X` ��   k4��8h-h6�g7m�      �-  ;�����pm� ��� 	  �ަ�I�X���Z�6�H ۰ 6� [��"Gl-�U* UU*�*�   8m-��X��M�`l�  V�*W����Y�j��c���tR�mPR�L��l�ɀ�I��lr�$k�-� p �``U�v��R���ˋ�6HE��( p  ���   m mi?o�TU_�,DU^�֗����^"�C*��(,�(
aO� ��|��?�|I�H��� �J=��6��vp ^�`t� ��hK� O�G�蒆@硡QG�	T� q ��HT8ShB�4�����ŉ��S�7�UC�z�x�� z*�8z>�;BsH��{�0�=�4�"&) � �tz
�G�b<N��TM�)�
���\��A�}�_0� �d&�)H�Q��h`�it.��G���)�*;⁈���	���2&�0#�`�'���U�@�H���*� ��|N�8���8 x�)�.�C 0�b� ��Љ /=@�aM�p�BM�/~�0���; =C�@y�M/[�= �`�H����!�<C�J �>� l��#`�B��OBqF�Ou�@���s���(���> o;A8����G�>"x)�Ђ@�>q���������'���?����G�͊�RI%A��
(�?�LV�B�D�)��(B� Q(a"CJҴ$�H��5��{����i��v�w�E� ��B�L���ŷ\ki���=�:�����R6gj�V��^bٙ6�-�v��6lգ�봵){[(�ζ�wf:�"�Nۮ��%��;j��GD�KɁ�ȳ��a��m��Ic��m�P�@���UW\�T�㇮�%�b��I��+3�2!#�g�s�m�{Aƣf����zòㇳ�mְ�Ue�m�Jr��%u�d�k��Ҭ��Z�vn��u�;3���"ѝ��Mc�Tm�3�mַR�5���Qh85Yi$��M�4��*��A4��+��3�"Ƥ��e:+�f{n�J��v2����m(�\�y��&��:���'h����u"ebƎvKE�;���J��V�U��j��t���*����D�\T�ٳ�Ѷі���	Z�˰Ҍ�$�F�܊:�j��Ńe"�; \�!�Ռ(���J���u����� r7UZ��^	�%CM���9l�Õj�O`����l��ʷh4t"��6�j:�l�۠�p��kG>tHU��	��E��Y;��oc[���i����<́�=֍��ԵUԬ�\��J�D��g�(8	��]D�V�A`�ph���wb���[�X15���rѳ�1[AK�[S� V��in� nf��-: �`YSW"v��pcqێݥ��L{9Ō��b��Wx��cX�=<�j��%@`��m��̑ۮ//����̇Z�s�f5�i���n�A*�@T����锣� ��6�UU[Pp�U�
��$�����޳TdCi�Yif�4���
[��8Kej�C�hP*tURYFUBeU���P;k�**�����S�J�M���W��;Z�o6^������ u��n�w	�mT<m�^�:��IspH�V�R�u�J�]M�\콺L�nכ	5��a��(.���
���4�*�@J��V��L��0�����C���N�*��j� �X�������pAA?�8Z �T"V�P���/|ؘ
'���j�`�'��POTty����ލ�Z�V�L��Tس�%�e������WnU�k�������`��۶�O����M�;`��fB�v�;S�ku�Q��{95YYG��6�gn̂<e�C6�$e�ч6M�hM*F���nH�b��&��E�p�',�� ��w��̭npT+�g�vU�CtKTXu�Y�� Nܧl��y��H{v*��-�ۚ�q�:�M�Qww�ݽ��0��;gv�>w*� D�FplA��Q@�H�"@S�Vs}���y�����y�r�u�J���ն��w-`}ݙ�R�T�I�w�`�o� ｸ��<���hr;�N����ŀw}z`����ـsP�m�۸��ڒ]���� ｸ�>����q`�&+���ݸ�ܖ��ۋ ����9��Xv{^�my�T\��e��mg���3��D����X�cݮ��==����e=��p�q�c�i��>����ŀwg���� s]l��v�Q4�����Œ���I���@�ڛ�޽�9W���U�y�0|жM���"�
Ik ��׀{��X��f��ŀsѶ4�Qq�݂��o ����>����� ��k�5�l�mD���w-�-`����������x��ŀy{ڣ�-���=�uǵ��;���u���N�E�cP�mgQx��8�{Y��
T!G�9���zn�����;��x<���lN��ww	%��9��{ۋ 淋���X�Ɋ�˂�X�%�%�*��=�ʺ���r8S0��.�FĔ�S��eB �Z�i�9��޸r�=�~����qkjՎ������swq`�L����k��{e�Wi�� ����9�^���ŀs��0	UK�h�+`%m�N�Ք��l��D��/in�mƼ��X#��ː���W5%��Ik�w���ŀs��0wvV���mP�
`�0{݋ �}z`��X;�ŀk�ٶډ�i�j�۬~�� ����7�vV�{����]qi��v�m��{��ʺ��xr�<�����?��8 8(��^�]�r�{*�aI�t�v]�u�o����e`��L��� ����/{q�����j+�����K�V����9��.��*��r�\Zv<�q��7H��nʺ��E���@�镀o�|`��R��j��+ =%#��LV�v� ߼��7����ό��b�k��z�Gi�q�;� ����9�^���ŀs��0|Ѥ��F6Gl������;�n,���s۸�lm�?-V@w`�ـw��X�w۟��ذwצ��!$� G�p�p�q@Ԩ�$\л�`A�C H`X)��Ҍ��j�L?����#Qq�St�,��sA���4X��z�=�8��{jW����-�G9��#��ll�+�ͮ����x}u���[<q+�.��y���
������uv{Z���]�Њv+�1m��nۍ�57'tvϭC��hr��5�^G�J�8z��q�IpnP�׸*�&��6��ι9^z�6�Q�f8��:�wi���v0��@�W2�M��;�&�e�x�T�C��g�+��c�����C���J&L)�ź��{��t�M{ط�QX�,g|����+ ߼��>��+ =���[��$w.�]�=��?U&��o� �t��7�>0���wI�t�N�[u�o�|`{ݕ�o�|`�|`���64�c�K-�0>��$$��6�������� {���]r���ݺ�7�ܰ�>0�{� ｸ��ݿ���7jAZ�݈���]7n#�]m�s�9ۮl�r[=v9�[�<lve���뫱�m]�;�Rm����� ｸ�zn� �4i&��������W~y����(;sa��TJ�a��ŀw�u��ޘ66��WU�I��Ҷ�����=��,}�L ��o ׫f�j'wn���	UK��X�0��<�{����_5I����}ό~�����~ŀ{�u�����Bjj%��@m�8�cj�D�m��흺��sJ�j�f->�6��j[����rK0��}�ŀ{�u��u��&+Nli�m�[�`��Y*��;�"�$�� ����<�����Y%�ܵ�{�u���R���-��^UJ��.��7۸���T�˱�v�]��5��0�L{�ŀ{�u���I5[��Gl%�s ����7��X�7^��ـw�o\L�b��n��,��J�r��ۄ���ku�W	�|k������F��.\�X;� ��q`��x��f��� �����`�n��i�۬�_r���~���K�=9� ��ed�Ix��T1����j��$�� ����7}��vn��@z�lR��ww�kUR��'L��_r�U������y+כ� ��1ZscMKn�,�,�7}��zn�v{^�z��7�g��u�]�;�^۫�6Uݭ��	7���g�:�Ç5wY�\n<�F��#L��9����x}�� ����-Rk-[�&����7g��˥RJ��R�IH{r�0�߱`��x�h�MV�cQ�jK���צ��ŀs�u����lm���%�V��9���zn�ޞ׀w޽0�-�m��ܹ�wq�X=7^�Ok�;�^�7w��(J�$�R���>u|�ݪ�c�49���=^�&z7�ykl��n��3ɋ\�g%�F�5�u��� ��s�G�GM������ �:+�B2�Z���\�;���b)���~|_u�L��g˻���0��2�@�.mrq�]�ԻpU��I�z8��!�.e3�{rܴH�@�`��fL�ܕ��pN^,c�+v�;􉑸r�[u0[FBix����ܳ�e7Ι���:ݹ{�n9XX�romck���C6��O[ʹ5��k=��ֶ��?����{ό{�+ �_r�7��s*�v��)+o ���{�+ �M׀���wɊ�ۑHX��wk�^fv:�sM�#���{�t?j�8����.]�X�7^ s���;���{ۋ :h�I��w#Q��X��<W��^�mhwL�޾ׁ��A�Z]��!v2��ݛ� ��ҷJ�����g;U۞��x^�N�Z��q-
˻���w=��n�\]׿:��m���
��.+/�����uHIВE+�O�s�^�����ۋǖͶ��-ˎ�wm�K=��^;��{ۋ�����9�,���˷%���l�{۸���K���.u�-VKw��%�罻��T����o��x�W�UIw���\��;hئ8���;v��ロ�]������ciu;����������H+w	e˾.��Z^�qx�W7۸�{T)ŭ(�9r�Z�}�쟿~8�K���2��Υ���"���7le������o�s��:IВ��
T�v��7��1�W��'7ѵC`I[�vm�=<:�E)�yD0>D�'�1��`�"c��$�.Ƃ�T���g
��*�����..���)&Aфk5Kr�̚h����jMY�aR���TB��{���!�x��(cRa�Չ�I��DR���ѭk+���Af `������h�� �z�p�Q�(���"�#�u�� ҋR����R���8�H)w~߱WT���GğX�cQ��[��\R�({�߾��)Jw��p�4�'~����(?2��~��)JR����ϓ�����nfb�H*�~߸qJR��}��R����k�R�=���pz��?  {��c?k7��Z��޳��);��v��m�W:Br��)�]v�6�h.�۷+��AFe��A���������~���R��<��qJR��}��R�T����*�U ��^��>e������o�ԥ)�y�����J>���R�����ÊR�����pz��;����)n⻻�$��H*�*���pz��;�߸qJR��}��R���o�*�U ���f��v)n�/^s�ԥ)���ÊR�����pz��=�=�\R��� ;	E"D���&!�	3��t�}�e��b�H*��|��>��Gd���┥'~����(		��~�/~��ؕW7�uJ��&Q�$���ȥ�;�q[�k�Ϸ�a��e��G��r�IK�����ћ]��f�Fo{��)J{�{���)C߾���JS����R����~��ԥU#~h����j;MKws*�U U���=JR����┥'~����)�g��9	s�ϵ��=	"��1]��9��R���߹�)JN���=JR�y�~�)JP��}��R��=>���v�n;v��ʤH)ww�W
��y�~�)JP��}��R���~������ܟH��e�r�˗��U �>�^��R���Ͼ��ԥ)����)@�}�}��R��O�t{�O!�}��f�����gg�TP�u�n8�:m�J=�e�l��l�����4z]vr���m�@z�>|}��3�L�S��6:�ݷ@�kn�s1�r�����װ] �d޻n�U��̠s�6�wd��5;�:��`�7ks�l�q���c�[�*���:��^"n�H�]3�@�	�^�2+���;�e��ܷFs��gUei�e淔qg�,��Q�[v�I��#���z�h=���םhK��Z4�96:�7 ��c���OU8F>�����ߞ����ԥ)���ÊR��{��pz����ﾙT��-�5K�H+w	y�s���)Jy�p┥'�����)N�Ͼ��(~����)J{�|j�E�E�;�]��YT��/�~�p�T�y��k�R�?y��pz��<�߸q�H)}�>�7p��d�N��W
�Jw�}���)C��}��JS�=���)>�߾��)J^��}��۷�V�N���R�?y��pz��;�߸qJR�����R��y�k�R��w������$�[kvӰ[m��S�n�x,�X�6-���wN���o� m|��1���z����R���~��)JO���=JR������)C��߿pz��?g���mݲ[�ݫ�r�U �AK�n�����'��M��Os��k�R�?����R��~{�)�1JO==����֍n�\n�˗x��R
��~�T������=H~���߿p�t��)I��~�\*�U/h#�'�)nEww��%)C��}��JS�=���)>�߾��)J]���┥'��e�}��5��f������ԥ)ߞ�ÊR��{��pz��.����JR��>��R����7�~�ʋ���l�.�LyCon�n�*��{��;N3��;��6�8+�nz{[��k{����R��{��pz��.����JR��>��R��~{�)JR}��7�ĵ%���!wx��R
�w���R�(}����)Jw�p┥'�{�ث�R
�o�?��Yr���.�R�>���pz��;�߸qJ{4Q#Rqt)�:����R��=���R
�
����o�r�\W�5�pz��;�߸qJR��}��R��ߞ��)JP���}��R��>=���Wj[�n��9k*�U ����b�H~  �=����)C��߿pz��;�~ŕH*�R�C� ږ]�����\m����M�����Iݳ��ԫ�S�۵v����nYqݫ�ܲ�U©R;����>���pz��;�߸pB����~�p�AT��F��F����ww�J���Ͼ���Jw�p┥'�{���)N��~� R����=2�vkz��7���5�o��)N���R����~��Ԉ-)�{��┥~���H*��@�Q�D+#�K��k*�RT���~��ԥ)ߺ��┥�}���(<TNAE(�1D40+E0��2�kP���o�@����┥'�y9��kf��̭�o{��)Jw��8�)J���}��R���~��)JO>��=JW�ߝ�?}��Q�����{��!��ݬ�{����n�m��w���29x������o���fV�Q���R�?{���R��~��)JRy��}�:��=�=�\R*�*��m5��aq^\����R;��qZR�Ͻ��R��ߞ��(�s<��r�G���>���*��*���kg�)<�߾��)J]�������~�����)O>��)JRw���ϋ�Yaq�v���\*�*���^RR�>���pz��;�߸qJ��w�W
�K|7��R��ww��%)C��}��J�I��~�┥'�����ԥ)w�o�R�� zG~���481gt�f�/Ay�VT����1�y�G_��w�|�l�$G�׎Νv�-j8U��nS��2��-�<�f^.�i�������m�o,ӭrhs��9Lr�v���׉�����7-���i�t��o�5ș%Yd���-��0�ύ��3���4�L�8kjz��θ�Ԉ,�sW��R[$���ov� ���_F����뭄e:Sw}���|N�̧nN{�ی�u>ջ�Ӡ7nLzɅ�۶�ۮ}�Hz�q�;q��v~|�|�����s|�8>@}9)�{��qJR��}��R��߾��JP���}��R��<L_@���I,����R
_n��*���$�����~��({���R��~��JR}�ә�ֶk[�0ު���R��߾��)JP���}��R���~��)JO���=JR�~؄��Ԉe�L�K��AT�W���z��;�߸qJR�Ͻ��R���߯*�U U���k~+��⼹/8=JR����8�)I�����JR��~��(~����)Jw��լހ��u��g�#ɬ8������](n��Hͷ%�]��n2v�v��j�[�e��ԥ'�����)K�=�|R���Ͼ��ԥ)���ÊR���y}��Y�[��v9x��R
����ė�*�];���04+�Wj����%(~��y��R�����)JO>�︫�R
�� ���(K���]̪@��}���)N���R�ʤI翿~��)J}���\R����=2�v]Ʈ
ݲ�/31W
�K�oز�R$�Ͼ��ԥ)����'� �}����JR��G�W�'z�kZݽ�g�)<�߾��)J{��8�)C�}��JS�����)<��u���ٛ7\���k֫����ݹ���ou�[��ػ�kj7�ٜ';�ٸ����*�����iOs�~��(}����)Jw��p┥'�{���)K�������f͙f�[��(}����� $2S��~��)JO}���JS��ߵ�"��n��}� ����y��U S�����)<�߾��!��}DvrS3�}�)JP������R���s�f%��I-\	-eR
�����*�T����ߵ�)J|��=JR����8�U ��/?�nՄ��ڷ/p�AI�y��┥�}���)N���R����~��ԥ)�ѯ��i����ʕ�k�b7hE�kۏm6��ힶ�u������%�qB;-��%�ʤH}���ԥ)���ÊR��{��pz���G��P~�A���R%��즚c���JS�����)>�߾��)J^���┥�}���)K�
>�}��Q�k7oz��)JO���=JR��{���)C��}��JS�����);��s>�����ލdZ����R���߷�)J���=JR����8�	� "HBI	���	"*B$�H$����Š�F�a%���(J��1�$� ������T��gث�R
�i��\R6�����)C�}��JS�����)>�߾��)J{�{���)I�g���3f�&�9�nkm�k�WccvӷT��5�uu=V{V�/[>���l����o�9�R���~��)JO>��=JR�����rR��~���R�������r�w$�����R
^�~�p_����O�߿k�R�?{���R��s�V~�A�������һm0c�v��R����k�R�?y��pz��*�)��p┥'�����ԥ)�-��������eR
�
��}�*�)���ÊR��}��pz����8�{�@s����UU(���J�k���JS�����):��~��)J{�{���)C�~���JSG\{bHRB�d�Bp�l�	=�)H^��a�T�<�^h
�4��*p�0\�$:GV1�a!N�R���d��HX�$���JJ�Id)� >�4�Hb��>x�1i�HH	J:֭a�l�����lH4"�	]%��D��Wr���ti� ��҄�!4����4bN4�	DE��,��IBSJAPPD�8@H��0�,I	D1K=fL��`-�c��j1	�R�<����z�1��20B�kXBB��Ů���@A�%�S��!����j.�u"ahp4Fh��1D�X�x:�BH����E-�;֎���&y�M��Q���;�0q�!'������5�,7�5b��5�)P�I!B�L���6N��B$0��5����HA*�3�#!qj]q���!K2��31�	$w��l��$@�̉PZD� �Ц�!�Vde�〙MJ�d�
�H�
_�}�٭Z��o{�fh�l�`kYg�#\ԡPQ��i�J�q�fY��n�wm�j񯁣fG*o.�'O.p��:�)^-	�9Sa6cy<n�>[z9۟nx��v��'F�r<2&6G]���aѴL(v| �3�[�MHM���5R
�Ʃ^M�2�3@��6�nx�'0ѺHbd�g�w����.�˻=]���atܮ�܇:�-V�B.�B �g��ia�-V��]]��['��\;䛣0򽝸U{�5�ʻs��T��8���M[U�iQt�m��L$�nʰ��AƦ��KP�WY%vk��U��M�:�C͇ �J,�#�/8Ւ2�[�����ksa�;i��y� 5PRԦiVH籊�.�.3Z��;U,Vʤ�t�PV�2JN�R`����.%�s���|�QCaZr,�<0���ê-M���!��՜��{�Iq�vŶ��\�[�"kkh����&�uO���aÌ���u�L;#���6!펐����.Mr�t�냳�zL��殧]����V��F�Sr��q9�v���^�Q���c۳4�����u��-��e��i[-3��M�����&U��9�a��wM0Kf���><��q5U5Q�h��L5C�ŤvM$���H�yT-�tC\�>�ʝ-I-ˑr�Ue{;��6Gi�׋�VW$����u�mv��ׯ$U�u��W[�ƙ6���m��ֶ���A설t�\U���X;M�R�l0l�jē��6�ZU�s�@�.��U-�U�kf���v�mI�+6���[#*�;����mÄ*ҭ��U�f�4���p&��W�@��e{�vn�0b^��*� e�����{�t��m�mQ~����wM�9|�&N�z�ں�a�M�2��1[oj$��Rv����*�V0��̽�v�]�d6G�b6�j 84m��@HO^�킔�T�>]���VPU^�y�c�'�.�>T�� R�����������@A[�C�N�y�h��c��PO8mT���}n�k{޵�EmCu��j�������ΩggGE��Y�����JR�+�͛����y��֥нѶ�q� �ƃ��o^����T�q�X�)c��#��m紬�,i��m��E���z;.�p9Z5�n8�n��1�c�A�ZS���;e�3�y�v�� �3r���d�3�6��R	T�Ush���n�lp��t�*:{u�a��c�;������-�M���;�ݹywn��)F�G�m��v�@c ��I�Bv�)�)�*�d�˹k�R
������JS��ߵ�)J;�߸=JR�ӦV~�A��ꞇ�-�mR�aE��=JR��{��� 3��?�����JS��~��)JN��߸=JR�w�4��\R6���ʤHow~�\��;�߸qJ�w�߿pz���<{]�� �B9��BA��j
Z7�k[��JS��~��)JN��߸=JR����)JP�ߞ���R����m�|�Gj�.ZʤH)s�oث�����k�R�>��pz��;�߱eR
��uT�7�K��n�T��{��q�(��,��m��ˠ��N�l�=���pT�Bܹ.K�\*�U-~ߦU �@�{�_����t��6{����wVZ���]�_}��Ȓ��I%�$�$a(��ZWN� ��Ͼ��>x����{��Hq��T҉CM�Ǐ@�����>��/t��ޑ����tScWj�n�`Ot���@�����s����o��[���Ht���������G�}:e`N��~��R�~�v5e������� 4��hIF���U����3�9�;�]�-�+.���T7@��x^������<�{Ȉ� �=��nj5j�t�.���镕@};�����_wG����!]�+Uwwi��t�����O���pU�ŝ��+ ���������i�{��UJ_O��"���@�t���������q'#���]�ϾـjT������I�/t�k��S(�I4:T���]��۳���T�޹��d����:��ݻ7m�5N�!�ݵV��&��c�>�2���t^�x/���'�#"�tSc���n�`��t^�x����N�Y@OC�RZchHvi��9{��_wG�N� �N���.���TU*SS�Փ�����������0�31 ���M�F"E�{���hHը$U@T�Ofk�@>���7@�}��K�$�Ϸy���n�2R:���=�m�W:K��.v��<v7X��v�+��,'*�V�o ߺM�9{��z���@>�=^	;�Յ�����>���~�z�tx��n��(�q'vU�4ݖ�k ��wG�}�M�>����J-ۺ�n��2�������k�ޟc�=8�J��QS2M%5U�/�n���:z�d��uUߞ��U�"���`��N�Fb���{��]��=��q��K�%l��͑��[\��I!����
�m6e�zuls�Ѫ ����c)�R�ѳ&��9�S��r�yzȍ&'*
�綧�Gb\�Ȧ���N��	w�WC�u�#��)Zi#7��u���yՋ�;����FŧS��<n�AԹ��@Β��F�R�ZX���m�Ի/J�Uw�F�r޴����RM� ��%��$�e/Nq2��Mr�r+���%����pXv��z�쵺�ۈ�q�كi�����R�
�$*�UU~~�k�{'� �1��D\ ��۰��512�R�qT�������c��{�vޖ�@7܄��`;����{��>���z[]�8���)	�&d�S6ӷv��I7@��"�=��^�G��������n��v�ot�r,��I wtx�$��^��V�m3���s���m��Jn^�n��%�<\�F��^�[�K�-�(���OIz�tx�$��\� ��EJ�w ��r���N {�}y:���UV����}X�����ޟc���"!!��j�0EQS2M*���y�݁�Kk����� ��t�������ޖ�@�N76�7]^{���`�A3S)E*GM.��nl�q�t�t�r,z��®�R�v�[m�N��c�����`�S�j6[�8�ݷ\tF�쥘�BFe�X�(wM<o/@=��6���Kk�{'��%!7D̓*fiT�UW@�w{��9�D$y��������wG�OT����m���4��uȰ}~����]�}�I7@��WS�VU�4݅����^�w�<�;��D/m=]��F�ҩ�UTݰ�yz�����7@�_E�{����~��z/�P$��F\��h���p��J�ݹ.�`q`��0�N��s��gmX'@T�S0�
j�{^݁�k�{��s�� ��䤱�m$�tX���}��^�w�<~�7@!"��ۺ�J�h�;k ��� ߧM�>��`�!"KH����;˷�a��s��ǵ�>�{v�q�����9�R����UUs��������~��ԒI-;�m��t��:^�������Ȉ��&�@�D�4�������#���Z�:'ms�8��tH��qٱ��i1�^��U���,jݱ[��<������@;���M��Eu\��1��n�_wG�� �{���G�J��EF6���:�Z�Ǡ���~����%��@�n��= �I�REL�hV��Ej���	� ߸���:-���i��"�K�57���t�c���9Ȉ�6|i�hzNs���F���K�ɺݐ:�]pB�=s�s�M��pSF�ݬɺ�E�"�HЄGG�w��@�Q`�khN�P�4]��UN]�Wڂh�ն�Zt�A�	ɑz�`�ڇ�.捡�oh�S��F��tm�Ԉ����n�j�u¯a��ҝZ �9�v�s$Z�4�<ug��7N`%R��]+�Fn��`�J�;���zV�i$cm�F���?�v�F�\=v��y�Vw:6�Y��vb5���j�u��u����%3�pIGc,HtF��Nk����t�c��c����y	-"�cV��1��G�w{��{�M���FÔ��U*��Sm��m�t����/ �'G�zG�}�tujۻ�`����/ ��:���t68�ǿX�qZR��1��7x'I���x�&�����}���PD���f�����F��4���K݌.���.�s���0@�=z���ufҲݧV�M�g����I�n�{� I�f�ޠ��!����xx��"}�Q��9���}��7��@>� �uR],t6��t+M�{� I�f�@}�'I��)�i�T�E2� ��� ��<zI�Q�tx���H�i;*�f= �� W��&h/t�.������Y3��:�zl�<��i�l`^�](n�SRz̓���~q��;���g��T��IT�t�ݻ��s��n�#�U_ =���+���Ҷ���mݴ��/t�.��}�=$� ���pe�4��M�t�@>�6L|�LvAo�-&�S@,�#��:����;��M��i�iuPPy)ڡAS��:�)�ؓ��:�WK�'`&�&�)EH�l/b�u�b�|�f��Z!Hp0�5�a ޗ1;^s�C�����k�:��HP��  @y� ��@�{D�GI��OG�v�a� 0};@�<7�N"�� *���׾{�]U�{���^��H��ҫ��I��c��#�$�7@����"�G�w�#�4���&��x�M�=�����ޑ���R�����.�Z�����
r�-����>{�\�6�˜���݁vg	��/p2]�E$;m���?�I�}�:I��)�i؆�?'m`t��ޑ����{��`/��#���v0Uf'���H�	�M���%�/W@��v�)\Қ�J���J��I&���XRH�)~K�H���GFZ�����ݎ����XR7V�����n�|�Gf%)��3��z�96�ݡ��s�cƛA�m�x5ъ�p/[U��HD14L�E)��U+ �{���#�$�7���_E�z�ґQ�aWm'cZ�c����t��}���H��Ju�]ӻ�Ҷ�'I�޾� �wG�{��=�UB�&ӡ!ݫ�������"������	=&�ޑ�vӱ4~N��"y���@����7sv�zq���G9B��Ь�?�1�B.F d�LBDL�B]b���1HJ�$j�)��+� ���.�]�`2D�v���r5Oc\�8(j��a�OW;�����3���t#[W��v�x��vz�8�RM�x�C,hF��ڜ�|D<q�G��qtqM�@�h�h�gZy�:����B�q��W=���&��$s�;ts��#X]��n�q���,.�n�HQ	�D�@6�-�CyK���]�єY�eE�������#�l�7Q��=<ɑ�v�b��!�e�}��x�?6N]s���n�ss���0:���z��Oi������[sGwݫ&5��:u�uv�^ ��u��w`{Ӎt�c�WZD�n��v�6�M��I�7k���{��`N���tx�=��te�j�UJ�*��d�] o1���G"8 �n�@~{�`}�ȩh�IQJjII��N���x}�n�^��XT�R ��՗N��o�}� ~����޾� �N���%2��I����3^7� ��l:x�s�[�b�v���o[ϞͶ�"	v�%�)m�w�ow��=�����V�}�����l��pzo�ԕs��~������G�Wkr����7v���*�t��?'m`)��}� �M�>��X��Z)tIU��
�ŏ�ԗ�[��7@���
�W{���ZG\n��]����;�tz�, �wL��#�$�w�� W);�lN��z}�v����o��(�]���9ۺ�[up��9�|��v�,n��v�@�����t� ���t��{��Բ�J�V� };�h�������_E����u)���Wmo���#�;�tւDz�F$�Ep�p�I!P��S�^�_s9Uם�4�i)I�]�WV�v��t��{��`Ӻf����#�=�UQ\�ݿ¦�!����^ ~��t� ��<��7@��s.�[Wi�cb�U{q�3Ãlp�ۘWVn�]e��8e{eϑ�f}�];-�G�v� >��4�H����>=���̔Bz���QP�z�k��{��;�t��^ };�h�ҡIv��իc��x}�n�{�Ӻf�}�Q����-��*���y�'�@=��l�7]��^H���� ��[g�ڑ�-˂�����3@��H������/ ���d��\���f;��ۃ��	�	~�)/K:%�Ū�-��r3��f 1Y-BԖ��ɮ��>�u�3�n�/c��A��X $�l�3R�&�����7vs�}� �N���ty����UEr�m� uv�{�{��>S�= ���t����w)�h��)�m�UQ�����������������V�Z`��X�����������y���\����~�UqD܈�����������o#�ⱚ3�vu�[]`��6m�WLkE�#�M�b�n�۵ìe�ה��v�<<����iv�-��� l��U�71�]��vPv�c���Q�V�fE�9�Q�m�Z�ݺ���.�:�2�S��Ss���'dJ�RKqQLj<V'ێNԧ��n�x`�Qe7�D�|ӵ �fsez1Y.��!	�
z��G*�8�����ؙo�����ww|�F�ۏ����z�IH����n{{m��-�l�v��; &X�Z-RM�T'�d�H�[�m�������/ �N���txW�)(MۺE���ս�>^�}���ryk{V�{]>���Dr >�̉��I�[����)��}� �M�>^�xWӨ	L�V66[[���?UW�>�G�w�&�/t������X $�l$�J�TM%T��t��|�����3@>� ������m/N1n%��oomlt�m��[,��uN\���+��,����v/w���f�!����^ };�h�������7@=%�*�S��M4~wn���3qG�F>��߷��W]���uWy�k�U���])+n�0Ux�<� ���cwf��g�yk{V���M�2˵j��;o�W��7@�{��)�������<�]�ݻ�[i�7uv���o"=:���ǵ�3�n�%��b ��ݑ.&�[V@u�mѺ���֒c9ӝ�4u�=���;���|�xDƭ�bn���@>�G�w�&�/t������t�Vؙ��= ��W��}�n���K�>S�=?UPw�.��'m��i6���n���K��^�
H�b��#�p���o~Ǡ��&��IQue��@�D|��z�3X��]��DB~{�X��:�%(�EDT�O@�<�VW��tx}�n���K�'��t�\v[fU�t��A���:ݻv7v���2�ݱ�뎈�#�$��F+���v;��//�{��;�t��^����ҡIe�.��i����7���~�ys��Z�Հ}�u�=�'P*���U�tݽ�>^�x�wG��>�G�w�&�z�锝Ҵ��v�M���;��U]����^���u�t)�Dh�����8������W�}(%;V鍍�f�x��tx��ʪ��~��@�<�Vɨ1(�K#Kl�\2�sca�tqH�{r]��� �a�V=\��Һ`�!��j��M��w�M�>^�x���V�}� ��U)����Wj������;���������G! �\#gU$�*��3S�16���c��s�^6���{��дWF%m�:.�ř�C�����O�|���/c��r ��c��i��.ն4�v��:n���K�<��7�W~{��W���i=�nϸL�?ǘ��AH�)�Rվ k�+�q8��Ju��3��W:3|SÛ��F��@l��0���~Aء��}�"HH� � ����"Z	"!��@�^�r3���9��������٩��a��;()(a�b�ܻ��Dwl�Xs��1"����Zj����`�B� >&�F�ɉK�f-�1*q�ą6	*��5�
ldٚS� $%_�6Y� v�B�i;�HP�%"V����b^�:�3��I'��v��FK�R�ր��x�hb�h��`n�kՙ�m����'Ŵ�5��3Y�t�Ҁ�;���\D�W4
��k�m͆��F�uS��y�3�a^�aC��d_`:T+mcâ������eU�2�;96��V���԰Zu��JH�;v��vP�㮻�x�:;{���Ĉ]��u���D�b�"�yݞ���Ohb��{FʩsL�ڦ�0��:� 뭞�c;ig�j��8Hۭ�e�凫�;Ǹ;uW:
.��n�p�J:u=��6�&���� VMk�8,ݝ�KR���Q�9��ZU�Ynp�����+�^�_[�E;wcAúU�%��lzۮR�\���M7�+r�18j�����P4pld���-WW��T8e�j��l�Y�C�s�j��N���i.$	k�x#�v�V(�'&L�����ϝ��.͝۞yCN�R��SN�"���B����)�E&j���kM�T[s��q����%���́r��ݺ9�p8��K�.%hVR�it�l�m�;�Y�T��E-�⇪���Ÿ� ��ۭ���`�'�Dx뷳�砋�ݝ;2ݖ�X+nXV��傕�;��;۝������t�\#��[��2� �����S���z��Q)<�lu2��'補k��J��)I�fW��2�<������� ��T�Q�[m���u�M��Zv�gp�
L�˻L
�v����h&���RV�:�K;=7,�m5T�[u�5��,X�� �9ր���3��lIub��R좼��:��A��Hy\��MH�j�X�����6�r�� �M��6��$ע��w2��LTʙ7)���Ŷ�D1K7d�Uݙ@e٢t+Ұ3�NCv;ˍ���l#��G+�	�����s��{g�:�gy�CdZ��VD-�����#lA��5�h�� �.����؀�T&��b�Tce���1\�b+g�y�w \��:��P�;���w>�������>��<����:��h�t	�4@<���z�S�f�:5�Y�{On*�������^9�B�Mәk����&ݞy{�(�x ՝��C��:m�oj� ��i�[q�iGm��P08�����gk��D�c[�;�m��r�+8{s�h�;q&٭֫r��)�ݣ0n9���F3�^�F��j�nLٮ�ݑn�U`<�f�jN� �������(+"�(�$슫$۲��vGO=�g�;|��7n��:�$�7Aό���b���|N蔧`; Y�,E���n�n���vշ>.��.�G�{��;��tx�S��HcMڱ7x��G�{��;��t��^��(%2��-����x��H��t�޾� ������V]:��m���޾� ����H�O*�қ�E�e���8�@�y���7]>m݁���+�:��ai:a�gs�mIƛ��$��X�N�K�f�iĮ0!��	�N�SJ�ŭ�X�n�|۽�s���t/T��?�[m:�b�ǠzG�~�p�C;��r9�"���v�8�@�y��b#��P(݉TL��)RUU]绷`{Ӎt,�u`y���bN�j�������.�?��I���tx��t�@s���HcV촛X�wG�_�����I�޾� �|��D�
5>�Ip�B]�-�e�$���]]�n]�繶t�SI�M9�W��L�!�_j�V���@�m݁���G.bm�X 6�KbJJ�IUUt���z�,˻�������T�Sbn�D�r�����<�w���J*E%�9ȅ�Eݓ�u�>x��(Q2�R�*eB��������`ǵ�/{�}���}R�IB���+�ř�@>�G�oI7@���`]������5�3�k:��H�>k=������n��������㓾?;v8�c&�7E�[�
��绷`}�ƺ�f:��������J�������z�,˻�X��]�w�H�@*uJ�*)MI)U.����`{t�s��K绷`{�,W�PFYn���I������]���N5�"&8DF�B��XCЀ�=tY�{���W�
�d��X�eӫi6��:n�����<����>�:��CǻS\AQP��TR.�1�[gA��P�m�VSZ3زq=��;Z7rl�g�d��<�v9bR7%�@�Ͽ<�}�������tE�*��һI�IM.���W��DD.r{�@�����_E�m/�hRP��ؕ�b�ʰ�����vs��8�@��c��j���[�n�����oN��}��.�G�UU{��$��+�J�������>��X�{������~� ��$�W��T�n},�[�p��).l�T��u]	�K�\A�WY-�ä�9��J�ڤ��rM�ӋY��,i��n=m��՛�bڞk�dc����Ԣ5c ��g2�s08���[ G<-�[�z�G^ã��΢܉W��nND�� �MY#�6�&�5uZ���Ůe�@�5�B|�ss�b��	Ƴ���������T;b�"�hݜS+=FK�Q��.���IT���(�-������s��v��h� nm�- f�q�mZ
lE-B�wq�����o�������zr9�|�^������I5TL�*�]�}�u��r!#�n��K��g���Dr8�P$�J��V�m�zt���~H�tx����=�ilRSM��`	U$��� ���������^݀6��.)9�I���߯�*J����9���z�,�꒕(쫱;
��]�v|��uy��=ct
�kq��e�];�\�λf�s�U�'�+t�$�1cǠ{��;��t�8��G9|��A�q�X�In�T�
R��[w.�o��9�I/�*�$�U��}��-<n��c����B�-�������{�yt���{��>�G�s�o���U����ۄ��I~<��= ���:n���K�%zJ�RZ�H�[�y� ������I{e�l,{= �{l�$�3\
�G(qՁ��ǻxqq�Ũ�r^P�����s�<��tt5jƕ�N���x��t��^ {��~��zG�{�]R���@��]��k��DG���}ď=ڻA��ۿ�#�"n�!mR���J%R+z�r�߾��:��߾�.��C�<V�WU~��=��>���}�II[ci)��v�����t����ƺ�,��Ձ�JKv���*Jj*i*���xۻ9�k�yfc� ���ۃ8�0?|�Չs��M�L���1��ƌs��ˉ����\v�ll��[vթao����.�@>�(�&�z�Ȩ�ɔ��J��M�3^�9ă��t��݁�e3��pA�p�5*fݴ�q�= ��� ޒn��s���������XҲ�մ�o ޒn�߾��^{�s��y(���.�������li7�+.���� �1��>�u�/w`y� �8�h��>3�pwT�ۭ ��lc��3�Bp�kP>���:�%�{N��Ͷ�_���h����M��>]���~�.�(Vݲ�щffh����M�>]�z�f:��r"8��F�)n�UUH�SQSIT�t��݁��s�b"��ڰt�x����?����Wot�����s�<�1Հ}�u��G"!|�w�� qQ;ɔ��UMT�,�u`o �r8���@����,�=!��A�&o�ϖF��G�[^K����=\��<���ƭ��t�6L��jzxX*{#8���vy�0u�e�=����v�FI5(h8�;
�5o`��.�n.ի>�9�Z���ֶ��4&.fH잎�!vQ��D1�ܷ���Vvɮ�}�u�콵�u�;�s�=��.v[.���x�B��kd�YS���D��:;f��s��N�U0�3f�e�n�o[�{�A������}o�����q!5Ь���<w�j�mW;[W�x1�,=�۳{p���V�n�,i���z�O�oI7@�wK��U@ywtzz�T�֬iYt��V��7���wG�ywtz�ty_�U�uJ6RU\S0I3Uv�c��噎��qy��绷`�`�UL���R�Jf��ywtz�tx��t
�_����>���%JV��j�1fc����7���wG�ywtzN�J꒨�ݤ�5vޮ/E̮�����m�Ϋ�B�6���F=b�۳j��QcB̷v����x��t��]�3o""#�����Z�����Kr_8�߯<�pIX��#�O\L 4 �����9���n��n�R<���M4�]��RO�wG�����t�����$
�t�mڵ���}��^<w`f:�lp����X 67�"���ED�SU]��c����9N��@>� ��H�r�Ҳ�U�zp��w]ctc���ܧ��K��6�����In�+{�^��2���H�$�� ��׀y��wG�oN���U)�4ݫ�wi���.�G��>� ޝ7@>� �_�����ڶ�1fc�������~��<QD�R�4����QE1�}w���&3a�l�i)�I�£��޺�oB�����u��sm�zs��$�#.htFU�pu���\�����PD���vP;L5.���M�܆I���p�eA�������hf����LX�A3О���F��\�:⚚ ��F��P:h���sG��X=
T�Q,#�s�����{���P�F/ IR�
�T�� zj��( �0ثꨤ���A��'���FOajrϾ�˽���B��ۻ��c������9Ð�z��&�z�{X������t�Hlnح����69�\������tǎ���q/|��Cx�;v�,�[x	v�V�n�Bs��Q{l����DC�~���������~�>]����$
�t�m5w���}��:n���t�?Pw�%:��Whum+m�Ӧ������3@>� �W������T"���G�������꫿}�|�<��C�S��Ug��Tz\�h�B�6ƛ����5v� {��4�����t�t���{��}�߯��~2�,��7^���k��k����R�����(�J�w1�������fg����Ӧ�.�x��L�'��6��blv�M�zt�+�˺^ {��4���	�J�:l�64�V�@����9w�=?~�������u����4�M]����r"��j�<��@��݁�s ����v��.�j���z�s����r9��߾�^���=���8����_��6.44�\�[���Юi���:$"�V���75����^Xݴ��E�tv�:P�r*�&���Y��O�O\�vza�U���Yg���ّ���\�JnSZ��Ƴtg�68��n�j���.5��d�j[�n��L����7l[�(֌Ys���wd��#i�']��Q��O��ƺ��
L���l����4�!K�K�Wi��m�5O{������z�w�7c�<���F��v.�뮣�r��зo���$7x���n�HY�LP�IR��Sʶ*����M��Ow����^˽��ӣ�=+����o��wot^�={lG#���t�^��DDqG95�A�UUR�J�*���<{V��]5/�^݀�=������'Q���MT(��{V""8{^�@��݁��/ ������VF��lM��J��6N��UUUW.�x.�G�I<�j!�����M��Ȩ�X��ͪ�..t[q�wD��;nݓtt������]sZ�����{�rE��������t���uWbi����w����쏚b�A�h�:QuZ�<wt���^��	R�lmmڷ��= �tx�t�?UU/t�.�G�OPJ��b��N���x������{=��:�9�A��]�<�(��&�Z�Z�{�r�K�"�tz���	��ޒ��X��t+��S���J�s�n�S��4{v�����p/3���&C���E�I;�x]�@>� �x��X��z�>�%��i)�n�b�ǠN� �:n���/ ������;�D.6�ձ:n�J��6N��r�K�O�_�9vtz�����ʴ�I���I��?W/t��{���G�l�7@� u:�˱4�؋n�]�@>�>�7@�~����Ѧ�	"j/�%����(�2v5������dM��vЛP��5W��~G���ޓR1����[� {�<}:n���/ ������)t2�C�i6�>x�����@k=��玻�Ȏ$fƹ�[TRU\�	I3W`5�g�5��Z~��ӣ�'Ӧ�����۲��;�xR���}:<}:n�~�_�y��xo����mG�_��W���ujE�����3�}:< ����N��r�K�"�tz��ZJ��NwUwH����И9�m�O��ݨ�4���w�v��h�����))����IMU��׷`b�9�g���G ��s�k��X4���*�i��7�/t�.�G�M������jK�Q*�m|E��L�	�(OՀ}�4^{.�՘�|��Zt�um�v��c��� �N���W�.�G�OP\���)ةմ���O�M�� �����G�(�RK~տ+�6H��v؝�KM�ؗJP9R���ú�!�t�^�GE3�d�5�,�N���A�^�N7�g.�{L�ݰ���;m���3X��y�5A��+-^�mXzήv�et��֝�5�6�����A�ߝk�]6ĵFv��B�"�Wp���Z�G ��p�,l�;�:�3�pL�('l���tQÞ6;bV��3Wm��Dٮj��C^�5���}{����o]qҝT�o;�l��1��/n�.%�L�,�Ol�f��d�8�o��������RL�y�� ����ӣ�'Ӧ�����m���Hwn����}:<}:n�w�<����}:�/��$��4�Y��������ԇ�k�jx���P��Jh��SI*��lG#�qo���c��g�� �txNJ��V�LLi��9{��w�= �tx�t�B�>�|���Sh܉�m��7n��n�@���m�`,PF�V�
o)P�,���t�e��n����}:<}:n�w�<��U�������}$y��}_�����9�� �G�E���	��%
)Պ�[I��	�����������X��t|�� uQU\�	E5vȈ��9�=����ڰ�:���tr�.S`��;�;�x]�u`ls���8��k�o���{t/-�4���	�i��Q.��ˠ���C՘�����;Aˋ��^w=�������"t�<z���	��/t�.�G�w�iF5vҷN�I��O�MҪ�UP� ����ӣ�:rK��E���V&4��{��"�tz?���P��@�ց ��k��.�Y��*$�@&& 8
&�Ę��B		T{x���O��M�k�� ���x�R���[i�V��������X��t��v/c������m�m�{o1�ӣ�?��~�Ԣ"""7��� �=���{X�ى��]��[��hޱ���q�5Q�$tX6������a���v�u�_X���^�=��:���9��]�JD_��6�5IS.������_�Հ|��@<w{��BA�C'b�*i4�����O�I~���'Ӧ����H��."t��N�ŏ�}$x�t��t�~�UV��߄�*��������|�F��ܖ����}:n�˺^{���� �+�W�T�eڶ�N��e5M2�l⣮�ۃ����竑É���u�^�rX�oZLLi��9wK�"�tz�����U@O�M�=�����E�x]�@>�<}:n�˺^U~�@}:���i����o1��G�O�M�9wK�"�tz��,T��Nj�ž׿X7���c���r�v�{x�\6fg��.Q3W`b�s��c� ����x������p�.G"s��qu!��0N�4l/H}�Ht�қ�:�{�f˿4Ȟ��#CLi@4��]�5�:І!�u. �m	��)��l\��pNK!�4�T�Jٜ,
�e�5�X8���xiSB�)���K=�A�FAI�z)��,R �(
��(�	�)����Z>��C#0�H8�R�cT%;:��;W"��# �	�Ĥ�!η��`�%d��t�0�JQ�%�i�Q5J�>D.;�wm��v@�(-�� Zl-�V����ݭ�u�v{7(��u�09A� ͻ-��m�u�D�l٫Dd���t ����`;8�(E��Fڶ�8�w���ڈ���Ni�Ul���U@\pG9jDgau�UՋZqW��n��#�/\2�S�.�E#N0ɖЧ��umٸ��)��;�k,7m�&C]D�v�<����-�\sש�g�O5J�`�w$��4�w`]97 nt]:
�����f]�8���-r�(��Eզu|�DuK��iI]�9�Қ`n�5ѷ���A��4�n�UX���9z��M�&۶��ѧd��nB%U�g��<D�=e���ݪ6�rv, �V�m]r�B��hVU1��UtJ�\Q) �t@ʵV�)D� �R�PDNm�V(IN�ToR��DO&1�� �e�v���)���Y��ƣ�cv�4UZ��F^E��4VvNȘ�*�;fw��\��)ɽu���\m��+�OZ;< ] V�e<b��Ҵ+4�ca6��ru3Z���N�Xzq��g�;��4��3ӽh���e���,�ey�m���r�v���:�cK�-��RvD
�e���J�VI���1���1�y����rtFѶ7UZ��*�U��^Ss�L��	����MQE��ۻ;r^y����l���t��TvC�.e4�[�ݢ@-��������c�{z2l����mr�r[���ۋjoT��xz	�
WS*�R��֙7��Ռ����rV�F��e�  ��-\V��m�	�n��Ji+`i$�MВ�F���敩�iUV�%��Kh[F�$�M��m�N�ehY�3Ʃ���';�$UK���B쳠 �v]���j�7]��띶��d��'�CQ�.+]�%�b�;f6T�q�W��݀U���
���P�U���,�5s�&�0*��6�2���*�U��@UKӒ�*�&���On���r7Zݨv�k73�Z��**�����JaP�^�"�>��� /���=)���A5Ҁ��%J�j���u*�����˸�i�s�[��l�vḮ�n��q-�v2\��N[E�I����������m��-�c�k)�.h��E������W<�,�D���-����k[<�N�s�ok�r�٥�+P)�ݯb;60:�#�����b��u�]�Ɯ��,�X�/-��H�A���[!3��]yx�:�f�� �;g����9�8���u��6��i�P�t1<p�g���}���񹜨oN�h�7��7j�8<YP��8q�D�9�c�=�-j�8w��X�4ݖ7V��w ��H����9�"#�17��#���L6l-؝*ŏ�}�<}:n���/ �������I)i\���M��Wm���t.�x]�@>��;�D��(�"��U�lr#��[���=� ���@�x��̀��J�AllE�x]�@>�>�7@�z��U�~)�v��-�!]S)Y�n0�h���m�ծƱ<b��:�m�!��Ͷ��m������}�<}:n�{�?�ZOՁ�:BZAD�QQ4������s��.*�UJ�Kۿ^��߯�t�(})~%���/΋��������}�<}:n�O*����vX�Zwv�{���G�O�M�(�tx��P�%$�i�۫�X����t�Dr7���1����{Y��w���~g����d�]�����ӧ��m��ՉG�Tڻk��s���nܫ����ITUM%SU`o����t����>��;���N��V[ot���w�= ��x�I�u*pi4Qi�j�����= ��xW����( 	%���FR@}M ��PgL�C���}7@'�xΠ:C��M۷��;�@}��@6��=�롱��ڰ7 'HKH(�
*&�UU�ͻ�wG�E����#�=��~�IYu'N]�91�nL���s�(ҳ�m�7㶢�qs�19i��$�i��K�pۿ^���V�7[ȎZ��݀n(�b��URX�Zwv�wG�t� �I7@=���u�!���bǏ@>��?�wf�#���{Vd���Jwv�tݴ���O���� ���ДU���U���dx��):t�b��ս�wG�E����#�'�M�=��Ү�(��&6����~M����z�ٺN�zҖ��F給C��^��st&�ce+m�wtz�H�	��k@=����1�m�n��Ǡcu��$o�v���fc�؈�P��	��
�TM$���o�v���]7��#���6��ٻ]�8M.'33�P�*	���s�f=�����`y��lDr ��׷`a&t�U2�T�T���g�Ձ����ݫ}��u^y���[�B:�qF?byo���\]l��BS���J�\vk]i�Cnm�<T	�y5MB�7:�]�qA��yv2��H���@�t��v��Ύ6b�Ö�zv8�n�{]����V�rkt��4m[�ۦ�yßtTuN�@��=�����gt�߻�8��Γ�۳�@p�a��%�� �Z�m�&ӝ\*��2E�����Ø9�q�Ua�2K�K�4�O��������ޢ�ĸ���G[����3a]v�Ǵ��Gn�q�^4;͹؀�NQ��o���R����`�������v k=��֒]q��M&�m+��	��������}�<�w��[L�-�v�@=��ޑ�����x��n�� �e4�(-��+m�����=���ݻ��َ�y Hj�m۶�[�z�H���� �c����n��Ir��N�����������<Y���5��'h1��q�	s�덍�	�HR�
*&�UU`{sv�,�8/zG������R�~R�YMRulr��<�~���T��J�����{߯����M�
�U�rӻjҴդ���_t�@>�~��ޝ7@�r��u�m���AX�c��G�}��t.�x��#�;�$����i�ݴ���}��t
��_����_t�@>�+�J������UmXնQG>7j��]�x�Z�\��sSGS��m���H�ݶ����.�wj��]����G�t� ��&��&S
-7m"ꧠ|����s���Q�G!��tc{��t�}�Te5m6��w��=*�߾�*�Ͼ���� �I��8�Q������ֹWY�߾�U}�__��jԶ���UU*�G}��8�ߞ��#��G�{�J%�K�e0@+�{�� ����#�>�t������םr밵�0�.J�nz���YӪ���rt��۔%��S�J���>{����zN��ݵiZjӻ��^��}�<�wM�wG�r��KR�m�N�e�'�������_�{�� �tx���U$wZI7wi4�n�N��=�n�{�<W�G�t� ��)V�M��S*��6"#�#��X��@�cݫ ���㈀�{�r�K���)�ݔ$ݵJ�x��@>��{���t������d��"TLl��c�kmt��cw'n�Gp�n�sv�!Z�`���NҪT�H��2��ww.]̻̾�{���g�݀{1�@��n��Pm��;�o �M�wG�|�tz�H��U~��=����ڲ�$��v�@=�����#�;�t*F�ݵj��C�����@>��t��~��U��tx�˩KRҶ�N������}�<��7@�u����R�U�F��\Q�ܸ]�9��\���҇/iKt���i1"Z�8َ�����0��>F\��"����4mn��}rۥS�sO=����2eP���}�S���ܦ�p�^u.9D^��9uy�de�8y��Urk'��n�n��zÓ7A��O�7ki\�Ֆv+i�G%�mWL˞e�a�#Kvq�s.'�`��j��sAgg"�vEU��vVU�g3�bb�޻������W|v��6l�S֢�����������v�b��Y?�/ÍϾj9��vx�� �P���k��~}�~�>����|�tu�����t� ��)mZM�.�t���]����@>��wM��k�����aj�e	7m"۞������n�lG"s���۰1I�x�JU��[M�v��y�@>�@ϳ�Y�z����~��&d*HQRP�Ut�1݁��"9̖�z��O�t� ���`��M���un��q������2C��N���$Ҟs�%�p�+����*��whot����tz�H���n�C�IM�m�J��޵��u�{���\Ts�
`�	R��=;;����?cw`�uݎDs��l�����U*:��V�]>�wf�8���t����@���i�m;i]����~��� �;���G�t�[Cv��e�v�����5N�����t�qk�W�V�M��軵ۯ"l�-�{n���0CqÚ�<썶�4��uص����� cX���I��V��5N�����t� �tx�JT�ݶ��w��= ��xwI������=?~��'�$3���ub�cm��&�W����l�=���3F��4�]�ڞ�в�]�X �8(G9�᭫J`my�ٽ�K$T�.�õ�����)JIS��b��i��c�&��p�p �f�{�M�t���UG�|p|�� �PM����8��{��;��@$��	ޗ���n�b�m�{�<�$�@>��ߨ��7@!�c��J��wv��G�t� ����=��lFÌp�O4�P���m���7 ⶟k��c����[&ס�nucQ��+Y&H��e�W$X����~�w[� �c����ryn�Հܤ��j��J��*Jf��fcwz�c{]�wv����*��m]X��J��{�<�$�O�����xt�tp���USJ�WCc�����V�]1�v��&q��@�z �|����������j�>��j�q�������$�@��)�wN�hL��ZcHI�ѷ�1��M�U�!أ;\\���;=�m���ͪ�U�b��1+o �n�{�<�I�}�<w���.�0��T�{��u���B[��`{��3w`�R6��VZt�V� �G�t� �n���/ >��K�wJ���i��bo�_������M�<���RH��I(��M��N�Wm�ͻ�7��G"2q���wj�>�u�� S�*>�"y�"����8 mM��-(�0�R����Un}0��H9.2�r;V\Q�n��jwtO!�-՝���v�z�ۍ��]v�Q79��I/I��I�s4$�7b���߿�P�n��rnf�pջK�l��� �ݎ^�9��:��l������;e����)g/[O�:��$8�����훮K���'<� ��֎s6��笠��U���v�M�Y�b��H�U�+.۳��NBzV@�֭�x
�C��\:�i���vDA.��:-�]����{v��1���ќv��g��/Q��K8ڗe�n�r�@��Lɶ��>�u�r"#�f6��� e&�c�$ݴ����䗠zG�{Ӧ�^�xޔT��m�v��o/@>�u�=���""9��s�=����~��v$Q1T(�*���������O��=����zG�Ot��r��C�B����<��z�9�卷V�������8��(��[�]��1�)��7�t���:I�L�ŗ��I�Eg�s��Fnڵv��N���I�}���9��Xk߿L ��W�?H��Wp�%䙛꫿>�|���h (&
@%�S�0'�  r��}����^�t�@�ZIDFҷi����j�٘����9��G8�ɽڰf�t�4�]�T�I�)����Dr"2q���{�`y��fc����	7m!�x���}��y{���đU��t2����{��N��.7E�v:cnv�pu��@�������^�uU�YLvڷn�-�z��x{1݁��s��G-�^�X�N�
&*��P��t�c���BF,{=�v��7]�s��=�k�ԁS@�J��8��� >߷����JIP�U
ʮ�O u�o�ʾ��몯��߶�nڻ���&�� I:f�}�<I�t	�"���JZ�������-<��	�< ��U�t��`��7m���o�� ~v�5�zKS�l���g��uZ։�gl[�omnq�[\vQ�&5ZX��T�S5V�{v�mt��� y#�$(�%J1۵b��%ot	�"Ȉ� ��� x�t�������+M�BV� N�3@'H�	Ӧ��E�}�@uOΛvڷn��y���B�Dqkݮ���n�y-��s��X�I)��#���bH2B�0U�@�[�}��꯽A!��6��L�ěx���UTk��`�����{��%"JI�Iӌu��uF۷!�I��s�Vp��;oO�Y�Ϙ.���IR��T� ����v]�p��X�:f�N�������Ѻ��WwV�+�m`t�:G�zN��N� }+�.�[�]Ӥi�f�<n���vlG99F��] o_�h�h\�ƛcM;i]��N�7@y-��<x�a�kݮ��F��B����$��%5v�mt\��z�� k���_{��u�]��d�0��d��B���R}_}��5�T0�����f+'^v�"��Y2t��E�nM�.جS���oW>nւ8�+��v]�94�zx�d���h�^��@����\����֋ph��l�Q>�h��km��Svv���H����7���8��l�c7vݲ`�Ų<���7��l���Ȗ��J���K���	�E�F�v�)ٷ�F�c����/v�e��:��y2��˖
�.X�J��UT�;��wO�N��ۮ-C���͟n�l��� IӽiKv6�N������� &v앷S�eUM!)��ׯ� ��<���E�}(ꔁ�m�v�m������ <�w`<��@�>��S*�]�+�%m��&�RK�	��4�G�zt��.�wBT��m��۞�?<}����<����Ѻ���Վ�&ۼ ��3@;�x�I������'�[�6VݝGY�ݹ����v�����n�q�r{u�z��K`��>'N�ٖ�`�,��3@;�x�I�����W�	��4x�)J1�li�m+��OI�Զ��QVr�/ 7Ӧht� ��K�*M�i�wmot&��<���DD��t?7v�T�
�JUSI
jz�Ȅ�k����� ����ˮ9x�@wT��m[�{m�� ����t)%�y�큱�r@ܮ)�P*QP�EB���נ�ݞ�@��q�7$�J2�ӎԩ�	��$�Z��T���S4%5]77n��m�@3�} 1��H�{<����QP��j���ڠ}������<���s��'�㣻m�e�n�zt� �I�_H����b�J�2� ��o�wϺ�?o� =����R�q[��38�n��n��׳aq���Dr���%"�)MQ5%*%M�7v��x�w����J�����t�I��c�x�Ϯ����p��k����ڗ����q=�cg{$�q]EE3����'�����w�������9L���ܶ�w0}��pUUUI����9:M�<�K�>�(�R�i�ڷn��y�z8`:M�<�K��t�J	����R;��,���IQϷ�¼Ͻ�\���}��W�@�%�T~'���aNޝ��bV�T�J*���<�9�{1���:gC��n�d�����]��֘|��m�ӌ�l>63�N7[m��m�Z�+�E��!��ѥ9#MO@3ُ�y�:�n��r��r^ N�T�%][�]����fh�� ��n��$� �{ŢY,llm���[0�M�<���U��~���tp�'r�T�6��M۲�݁�۞�ff>����-���̂�)���&�+w���4��[m݁�۞�8Ϯ#��"�9���_Wu%"0:9���\���=�=6�JC �jl �e��OpS�a'{3j�H�	B�=��	�)��w(`�� 7��h�<2�Հ��;ؙ� 9�W�pX�4�D����؋�����j ���}8!�m@6��*�����~w�\�o{�{��y�x�t�����([C"��յ��rX��:W'ZhA�'h!I��q�MU����f�kJ�M�CV'��It�m�l��m`e_7b�:�¥Ӹ���6������!������x���� ]&ᚨ�ζ��[��s��j�2��tH�q֚i����;�7+�-On{6���km�5ێV�&�* �uYY(�nI���u�`�ܑ����fR�tm���+M8�;t�EE&H(��c��|lnB�8b��Τ��U���5���]e�iLBg���^�Ʀ���Xκ6Y�:|����F�m�]��B�{S���-�ݸ��6.�mv45ˊ�����Y�[<mD`�F$Uņ��9�j�$�*�X'���V�UT�&p��ĳӀZ��T-S���P������չm$�͍�,s�T��tB%eG!h�NL<�3���ԫ�OWF�W[n�"8T�m�p�m������̏m�m;�a�*�F�[+�7��
ڸ�θ1�U�!�tV��s�gі�-ۓ�0@<i��]bol�8�In��D�L]�=������U��E����Z�E���\�okw����m��	��i�I�l���UQ֣$�H V!6|�u.���kj���/b�C�PX�"�:��sp�d��V�Rړ!!��.1��K�1�s
�SC=�܈��<s���K��;B��ђ��{��%���[����8�ݭh�NՎ4�¦iݸj����Nkn��o�8�ץ�km��h ��A��g]��Ӟ��0 �l75x�ƴ&�W�$� *K^�Hen��թ��iIj���핥^����f���K'F��*�v4ܮ�W���(����D.�3 �;��c����l����[���i�m��zn1s����bb�y8��^vV� Ȁ�l�*��VÖ�����f�a�>�q6���ts/��UK�j�f ��E�ۡ`�Ssݳ�9k,�튧\]���*�����x��@�"���)�͂@��	�_OQ�3��t���u6e�ֳ7���@nJs��V^xݭ����3��[w4��>��1Oas�H��3��	��vѱ��/��VW�r���`8枈+��2u����b��Bm�[��t�E���=�;���q���U��Z��;	�vz��ێX� q5�]o�g�8˳l��<�'#V��6S4�.k��@5��Wud�<<۶��jJ��s�B�v��'�E5��;���?4w�"q��]���泎�PS�ܞ�#�u�9��	j�-�Z_7)8��I�#-bq��-˗2K�π��V��n�&��31��nX��D�J�L�&h��w��q#��@7��33��9�� �jى[<H��	�Uv-ݞ�ff>ټ�9	7��@�wv��p�S5H�$&*UT�=��`f:g@��݁�r9�۞�ju\�%]��Zy��wG�����w�Ż�������ozJ*��&̖�y�\�<\m�vS��-�yFh�b�7�}G�T�۴nwc&]:�j���[o���v�&��=��`f:g@o�ID�wr]��p���<�����H�Iz�R�������>�Ztx������Q/젷e	7m![� �'�h�� ��n��$��)ZM�i�km���W���0�&�RK��t��P:�.�1�һhv�gI������3@���Go���C�&ϝո�kormn�{$�,�tvǆJ��qѮw"�O�X�g`���m�۞�g�l�L��D ��݀<\�4�RI*��f������$7��@�^��m�:��.dq3H��EB�|�:��~��*��~����{�I����0Ţ�0gX�	�����('I3@��B��l�n�bV���Ȉ�"!}�v�ݭ:l$<o{`7��ސ�Ҧ���i�v]��=#���G��� �֝�7v���)7�L�v�N�v^��n4 S��H���\��/N� [�a��Bj�̢�\��� 7��4��l�7@��E�R���Ҫ�W5U������G��n���� w��h���\J��ui��0�&����{�f��0�Ә��J)(UUv�,�ێ�}��~�U{����i��\Q��	EJx� ��C�����U���֥�rH�v�wo 7ۿg Ku�:�n�9mt��P��4�\fƭmϳA���s���u���3�������l'
��c���)�7��fp߯� ��7@�� w��h����M���������o���q#6wW@7��;��~�;�T�ۻm7n˷������}�b9	7��@�^����R���v�J���t��8`:M�=.E�}�Q��M�i�km����< ���f��r, �wL�"K�\J�i�'�s�qF���c�v��ӯi�%�\���]t�6Ët@X��Sfu�*tI�ݤ�]�.�v۶PÄ��vU�vw�ً���V���j�vM�[	���e�j�kg�5��W6�XMWV����nܜ�W'	�[�����͠�gl����`�葻]�kX��+cH8^"�+OPyzy�[iVvض�st�0g>��:Iѭ�n�� ܜ��dL�%�/R��I5���+��X�vb'�� �v���:���k� 3[w<�m��{g�^��-�
�m�_���ϫ�[] �f>�9�@f7]�DBǋf'fxr���*���͝�� �f>�t� ��n�O/ܬ��I�B�J�k ;�&ht� �t��z\� �8��U����v%�7���<��n��-���AȄ<{��3%$���T��n�v���>�&��"��I��#�$%u��IF$��wg�ST�	v���<��ݹ���9ۛ��詭�&r:t�Rb�p;m7n˷��Ȱ��f�wH��I������m*�v�J���O�ք�$�~U�;�߷�|���~��PyI/ ���uJV�j�n��m�ht� ��n��$� �wL�=%�Et�CE��o�:M�<������#�>�E.�+(E5O�T�{`ycs��c�{��o�Ў?�/g}�+G���m�b����ugRݣ�\{(��<����� ���z��}�cu�-�w�E��-��jqd�I��[�,I�f�wH��&��"��t�޴��m1���RS5]�7v���o""xs�r#���bF0�2.HP&�ő{�Ԋ���>"�C�-��߹�s�0�ƕ:M�����v�@��ct΀g�ln��/ͻ�23���ˡݧm%v� ���h#���n��Ix�|zJ�N�&7wC����=uیm��tu���x�G�)һ���۰!��n�VR��V�v�[o3@���v�nv-����װ��j�TST�ـo���yt���t��0�U�e�T�N���<�9����ds�c�t�n��s&]�v;�M:I�w��t��0��M�c�9��3��%U�UI%�7��߈}>cwN��'y��{���$�ˤ� �wL�ߞ�{�>��<쉿%����#ն�࣬wl�ݷCy�[2mź8�z�]mq�G����	r�cj�7L�l�>���۠yt�����8`�ƕ:v�M���v�@��������:��ޤd6�g���;in��g�{��9�D���=���dz�R�SJ�i
f�X�L����=��t5c{zX�R-S
�"�EASG@�w`{'��}��~�à\eG9�`�W���T�u�H
ݿy���;q�viz:�%�F۹n{sj�W�����^-����)�h�ۈ������G.���uZ���K+l�2�S�`�vA/n���p;0m4bӀ7�s�B����&�'N���W�pdx6���=���n�s��铭;�ධ����+�����+��(��nt�)/V�\$Xva��xڞ�4ZN��e�vrt�����www^��I$��v��D��\j�ƭ��R�0��۝�W�w�z{�^�����Ʈa����B�SU����k�{1�:�+�~�w`y���w!r5����n��?�I$}���>���d�]�9 ZxK����Ҳ�J�yZ�0��n� ��e`���]��-�v��[07������r�t{)��+��иҧN�n�ݻ.����`~���#��g@��à_َ����į���P�2;�^=�Y�ƻ8�[�;iv����1�3���`v�����R`J?���Θ���}���>����QG�����ݻ�l���w��ƒ��T�I$��\DDDG>����]��[]�����*�TϾ�ˇ��,w	ar�����Y�z����/�Xt�	����l��[{�ywK�>�L�{���=��76geT�S*
����>�>�@�s���V��;�3'���w�8��4�%��ݹ��a.�cŵ����ӎ�y؏>��;r����+���ɹ��}#��{����`{�V�ZI�wcj�h`���#�t��t��7������N�ƕ:�۶�r�%�k��`���Ĕ��"��0�c�<pזQ��&2
�	"`�����e�"��1����{ۄ,�Oq�͖P!�����y�������sd��u�$�� �1�[�ɢ)�	$�P�VTj����%�n��(������"� �#�1�ʤ����+��Q@Oq���#a�V@L9d%"�Í'���9�zs�º{#GGbI���)
��m��o3�a����3^���W	n��k6��4h_@�͚h1����<WF�:�ک<;/��PY0�^!R	C�X�NE��i3���Ѫ�`�Di�zْpN�@� ��RBk�ktGg֖L1�pF0�&�l*����!�B�
����Ap�� h�8Ҁ&">����i*(/s/_zt��p!��C�N�E�OCa{�t��t�ٷa��{=Ҋ:����6�M�V��hH�T��}�g ׻��;���#�d� �߫���C�7x�!������Cwl���-=�/\c�Eؚ�L��ƭ��b�s�>�>��Z��t��Z��S�6Rt���9wK�>�L�{�������I������'��B�j'h�.`ǽ��y��@���v,�= xz���t��i*����0��M�;=��r����LJ?���e������ji"&bJJ��ZI�UJ�?r����g��&��Cl�>�����ܻ��zLX7oL~�$�H�N+p���v)�<�g�#��A�suڻvv��la�m��m��6��fiS�m��n�]���t��I��os� ��t��p!��C�N�Cnz�o�Ӝ������v/c��9�${`�\j"UR�USJT�Ł�u����z��}/ ��e`ޤ'ŗSAB��)M��/{�`4��@���:�o�����L�J�"�)��c�����t̬:�{����m���ゴgWm�����FzB��/7A�7\A��]�/J��j�u�^�ˮ�P��vrq�H��ݸƞtìu���BP�&�^M@ֱc-<V�g��w['m�V�%h_)u�	n.��g�ݞ�{oB����S=[��}�펁6�ľ��Q��8���јݑs�g.��vՀ�������fh����14n�΍�����ljz�a%+�k%>�4߾��|������Ӓ�J��]��Y�=�3�lu��s���h��`��,�v\@s�����<���,��{��/2��}���c��f���-]+.�_���>�� ��t��t��I��{֒G.e����0V�ｎ�Y�z~r#���w��>n��3zT��m���Wv�@��/ ��e`���>��7@�	҉�t;��[w�}�2��|`}r{~kQS�K�ڒ9lM[D�r��y��V����n�J���1i��v�=�%M���{Z�8`}r}�2��&;��R��dv��0���8�W�
?��t
|�uo:�Z�]y��:�Vy��T�!O�"�)���og�}���+����n�76g��t�EZ'v� ��e`���7�o���~�／�>�8��Zu$��>�� ߽�t]����+ �u>��s��%��Z���k�C�7
nΟ ��%�)ns����'�n׈� ��Ln�}��n���/ ��2��>0��*v6��e����^��e`�|`��n��8�T�wi�Hm�w�p�]{���`=B��`�1�ȎG��u���\��@�EU3E6�ݽ����r�K�>�L���B}j���-4ճ ����s�f��n�:���yf��TQ�Aѩ�;�p��\�4��H޲j玠q����X�&��<r<C�a��ԍ}}m�G���p�&V�������_��[���&������7���>��7@�z�]�Z�V]:���+@�s����/t��I��}�I*:���I�E0V���t^�xޓ+W��d�A�CǴU�D�;� �B�J��ڶ��V�@�}�2��>0��M�$��E�.���=VG[l��7�S�]�m ]Uǔ"����Ϟخ;ps���G]�&S�m�?; ��� ��t���^�����V&���ս����{������&V$N�D���]:be���`�۠r���}�e`w��)E`Я�wM��{�r���}�e`w���M���.�m$�X��5n��}� ����;�o����L.!U		XHVQh=�ϰ�f�k2��6oz3�A���(���z����
�gn.������rV�:�zh�d;%��q�ϩ�X���޹z�g����jb�ڜ�
�S���]����Y���{ 8峫t����)�#�.�y<]���.N�t�2X� tus���j3�q�j���4mO[����5�mPnby�-0�ZX�>�f��a��jNY�6�ϙ��8X%*��P85�Y�kz�!ꂇ��:|���0���61����m�lx#�V�"����l�V���[�7�Z0�,�Z����>���`{�7@�}�e`z�J������`����M�9{��t�X��IR�J��ڶ�v�v�@��s�>��?#��%��g@�c۰3�P�F�ӡݧm!�x�&V����������uwQ,�Ӷ6�j�ց���wM�9{���2�ԩUw������V�v�ƬM�v�ذu�Nڂ�ق��=`3V���ٶ�C#�9�
�R�,f=���@��o9�<�t{��f
B�T�LUL�U��}�|�lC�p%%��/>��9G������t�)j[T��]'CM��I��}�|`{�7@��/ 'z�]�+�����+��Ӝ0�r���}�e`�I*:���Bl)�l�>��n���^�I��}�|`��s����moPsrV7r�q�ݺmg:r�\&�]��D�G�M�W1ol��5��9zK�>�2��ό�{���N�n�Ю�m�x�L���� ���t�Ȱ��;��bi�l�/��{�����N�R����V�/����XOL���"��*t��M5l�=�t��r,�&V�y�OIJ*�I_�v�6�v�@�\� �I��}�|`��n�}Ԋ�B�HDMx��_X�״s۶y�)s��G��qvđ=Qu�{嶿,���I�J���� �I��}�|`��n���^ N�.��*��K�3ذ<���r31��'ut��������� ;WV��;�o�������!/=��@��g@�p��Q*jh����EM]��9�rDG���=��*��7����"��¼������˨WP��B�M�N��I2��ό��M�9zK�%T�ZU(Ҷ��&�9�wZq�n�Q���;��v85�5(i�ݫ� ���l�Ӷ6�j�ց���r��������X}�E>�®�T�R�4t{���9	f��n֝��a�č{��D�%<�TEUMT��f����:��à}�c� ��'*[M+��I��w�_�tp�>�>0�r���ޢ�ܱ]�Wt�U�Q`y�3�-�r#ُ}��T�+���_����EU���(������3�0W�7���ƅG� ".���@�@��������QEU���������7����޽�7�����e�������U���?��ʪUJ������g���?�EU�AQU���������?��b����o��/�ۇ��9����>����
�$ JJ$�D�-
�,��0�H�*$"����B�
��HJ� �
A
$B�,��*$ʉ"D�����(���BL�! R#B%�)H!@"�L0��D��BR҄BHI@@@J�#���!K0�2H�J�,�"�B@@� �� J�� ��!"@@J@@J�H�	 H���!@!H* P�$! J��!(���Q�@�BD$A�%� �P�I�(@�Ba� B� !	�dBB@�@�@�a�d�&�@�@�F	BB� 	�!�d@� �%U�a@�	�aHB	HBF�!T� F �aI��!�da!U�e@!I  �%QI@ �%�a �%�!��D�
 @��iFQ�$Q��!TQ�dBP�d@A�D%A��dQ�d@�`�	F$�aXF�`IF�daQ�Y$! a@A�T`Y @�a	PQ�FB!@aQ!��$	�	FA�$ �!@�eB! �	�aQ��	P$UB� 
�aAB!%Q$Q��!VQ� $!IFe@�B	�		@��d�I@�$$Y@�X@�B  aPP!P	@�Q�	`BEH@�$H�aRD(�H@�P$e����������=��]�������ӏ�O�|������d���f����_��������������TU_�QEU������(�����QUz#?���������5���^�|;:QU��?�� TU_�����GQ�?��0EU�]��
���}x����#3��r���������c��ˀ**����=��`}���O�~<�� ��������} �������������PVI��Z����V` �����]5��  
��� P 
 Q@ @T(��(R�P � 9QD�B���   ((@
�J�P   �      �   �� �� �   `R�DTU�"�T�>|\Ͻ^�<�_o���S��x���ݾ����W���w�-�C�O\���ΐ /��v�����`:(pۯ���O.6�����>�)W��������Ş�6��� P{�EP� H�� Š*�>�n��h  �� @��H*XP�p � � �  @    �  �� �(" �1  � � 9 �  � � � 0*��@H�����Gs(�	���5��}��Ϫ���P=��U�z�W�7��������}x� ����oW�\�� �{��m�3�ַ�E����o}��������:�����+�� x������5精�|/}�xi� ���B�UTI�c��$�����Y|�s��;v5� �%��J�g^l������}�[�
�}�_.3�V��� n�;��ﾻ��o�>������}��<v绝�wf�<����ӏ7ӫsuxޞOK���������)R�T))D� ��Z羚�N����9������}}+�w!��׽��z��������o��<v^  �x�KǷ��uw��^>�v{�^���N���'����
�o������J�e�rt�[�^   ��*m�*�  ���#jJT�  �=U)iF  '�T�4�(0� *�J=�R�  �!'�)$@��<SaBk�/�ԣ����9�K�SP��w�D(JB�����"��TU?����DU�uEV 
����y)���!,�ĉ	��"$j6	!��6m��Ed+I!$r?�s�1����"B	�ԃX:~�~��ky!
J~o��?��V	,*Eb1պ~��L9�_��������u&2�
����u���~����|���(H0
���mj ��	k����uqM�M�U�.�R"M�B�X@!A��f�����A/��M͖��j�/���K�_ξϷ�� �Dk��x�ɍu��)����
P�aB��sA�+���4BSS�K��1�4��Q�͖M�fBa��6m�0ѣ﷭j�"��Әv�f����&�(h^��n��$? �bh8:M��N�s�eϘm�t��Ò0I�Y"D�R �]��Ɂ��Dؑb$�E��du�jB��T�`b@+�l�Fiu�$f�dE �i�j��17����� �4�$i�����6���J i��y���~���	�H$a��nol��(biE����l'�2,�e0�0Ӵff�ٌa�u4`%��.�d�[ˌ�$x��3Z!����ٌM	��!��d$���fۈ�&Y��@�*��X��l��f��L U%5��2%�$��o0��q�a�)�(K�C|�񎝋���`F�����ٳ_�B\�3�c�q!BH��.h��.��١����[�E���rr��˴Ms3��(�=�dB������\49�s�\�0�ϲs�̷��:�B��AήE�emZ"�X@�S���̦���k�����&��Y��||Fe�0���J�-%11b2��d"Q��B�RHP�!\Ӹ�����I�sH��v�"Ɵ�f@�P�n�-�)Z�H`�P�%J�z�I�+��#�}�����&��n5�2>i��p�Һ�H>'��7߆\�K�iY�鐻�}��f���'��5]Sz*Ege�D�v���cEK��Q�*��y,���sy�j��L��d01�X��� �kX֬-)JϦ��HJ�����!H[ch��\4�AA���)�$J� ��@����0�����#$�`B�c�Ld��� ����(��B������t��-r6�k�5�BkI8D,jB�HSb�
f�1��:�S���X�n~��7L�.ϒsﻭ}�s����`c�J@�iCeqŔ�J�_�I�N����)$@�~�7���d
��"�.SU�_��;����>�	n�S�%���
��@1>�<�H�]�]#�#q!�@��D��v
bh�$�� D�2D, ��D܎Ԑ̏�G��8B2H�,	
�z��c�x����� ��Bg3:��/��1`��>�a��5����B����l�Mk��ޖ+�3��6�ن���MD�Gi
��F�>8@�C��y�)�������^N5��\�1�WPF$\8Ƹ���-U���EE$2�w����F]� ��5�w��YxR����6~���D��	�"W5�3#(��~,���6ZjZSi����)G�P���F�L>aLћ"P"T�|�VR�$4�vs�>aR$0�㳉��1(a�g��D�Nӂ|S4���"1!C���Y���B����z��h���
B��`B��F�E14�+|Mg	V�5$�in�iXr�uJ��1Ph#��ʸ@����������x]o9?�JB�6˚	u�$+�I��ވ��SE�����yN2�Y�V�pEn+1"Um�]��S]\�� I�8\e���� G�c "�JFB.:�w7��I��W�)�O� F&���>H8�����!Hi�տq��`�!u)�u��E�R"@�1?a\�4h`i�`XBR~iG ѳF��>��!.D�7�m]��n��D1D��I��%�%�\�$C���Q�]9�l.��5��XG4~�cP#P�SN�i����h?,����� ��x�`���k����>�b��8¤��B @�8�������r4!y+��3P�:a&�3�`HA�t���BRG!S	d"y
f�7[�:0���(B�||l۠�}:����"����qe��U�Q��W=��5���|�`|���Sm��F�$��_I���p6�0�k����J�rd�MpS�s�kX���.��5!�pӢ\d��0�l��]�cp0��~E�k/\$�0 F�&9�\��+�#��_�e�XP�1����)�q��|������!��.c))��Y��ؐ�}Mad�F�������Ė	ą(H�9ׅgm��$��/7"�
J��j�� C�����?��[	��v��]��#�������c�O��h��M&�������˭�1���p�QĔ�+p��)0�"B�.RTӎ��
��\�tm�M\&��&D����,�k�d��mZ��R7.����%�Zm�H���(m�Q������>8c ˘RP�D��%_���jB�2]�� �d���q:����o	p%��ѐ �#Á.j�>38|k�����;̎N�ڻ��I�O���d�I#c��8R^��:�cO�ۚM5L:(U�Z�*N�)[ΡM咲�F.Ga
`B	����d��]��H\p�,t�t����fϘ�HS�%�5����N ��[�o�C�����0�S�Ȱ#�)����q��
��W{<\y�m�sB�D�3��_�o>���J����aP�X��cX��H�R,!$��Xc)؄%l����+ŗvH@�R�H&1Y���V!e�rϷ8Œ<af�X�ɭ]�F����5���A�q�L�SN�}ro�L"D&���(`HR�b��kv!��D�|=t0�@���&a�0����R��FY �����	a� ���_�$�2A���Kahă!!�"8�9�u��ɖҳ�1�.XZa+�.��s%����$��
�Fl�����--���7���$	wi���k��oEm�}'��Vy�>��<R�MݮU�#Ev]%&A#Q	S�F�D��)����W@F"�"�c?�"5���1+M}�:�̤ \���q.2�Ʊ�*@���.�h!`�(D�D�%~���	�_ͤB3\�f���?O�JŠŀ�K�����!�������r�^C���Ӵ�\H D�)52G>&c.0�2!�L9��}Nr�5�٫���J�rs�/���.b��N�p��gߒ��uXSA'�k�a5!�5x@���,�����{��|��$�a$������l�,r?-��$#S�#)�ǁ)��0�7��d�Ll�PGH�PLRe��}��J�"�fBP�a����,�@)!e&0�!�P� "�]�$��+�|V�B)]�V�:g�����9���;�\!R4F�:HaM���$ne�㫎�bVP�G[���ə�d��.���%�h&�1I�eLt�ġ����v��ĉ��E^T
aT,B�WhU1#4
ġ���]&������eiƮ�<��#�;�̩\��Rɭ�e�3�|�$Y "�M"@����p8���Hd���
0�*FĢE�J�����/�6O�P�$�<k���%!.�l���tm��L.|[n���k|4kXr�s��z�u�����++H�!	�HR��XHҰ�B2��K-IBS#Њ�"	]}�5��4 �@���}�]�~��H!$8����7BI[���]���	YM�)���p�l+��I�{%�
���<xt�K���m��e�ӳA��bh��4��ѽB�X�0�љ�u�a��0�ϲ'�9���p#�q�H��ւ@�B��@�Aa5��j������\�5��Fo�}�CM�$.$������� 6�	        �8   [@  �a�      �  ��`I6� p      H ��� �   p      	m�  @    ���       m�    �0�tnE�� ul:�� r��l�l��gv������vbD��-��p8V���ۗeve��[lJ�1� -�!�lH ��` �b۲еnͤ��ܖ�x �9m^�f�IR�6ۜm�RiM�x�j�I�-�`��m����m���5kc��� m٫g��M�I۪��b����N�nb�^��diV�a��ٳm�j�3�q&�$:E�5�-� ��M���m��ph��BKrl�����e�5P孁˨�J�&��^m�m��䍗�
��:f�7k��n���ԭ��ۉ��e�o=V8瞜֭�n0������E�O=��E�Q��C��xm���λ+�{r�u�������2�V�gC��y}P�GjyV^s�.j��m���j����N�N��/��U_��)^�Djn��ny�m�nq�k�N�o^��n��6��8m��l۷�>��m�֮�"�NkwC I!��sg[mt.ȶ5�=f��]�ދ^r3g$K�Y+t��dt�\�"m��{]t[����i#���mzf ����[��ņ�.�����e�{%�[�É��.�nݵl�D[7��tV���-�A�D(�;�n3-�]��/sVqڞ�va�ո)��ʻ[USm�Ŵ��h��l�-�  �I������ n��$�h[�lݬ�$���8�h �t�ְ(�t����]nRsB�e^v���]muH�eUٕ �����-���k�MOlp�%f�kj�dm['I i� ��K���l��l�8Xf�I �:��`��mm��c��۶� 6ݜ�d $rG;l���N���f�qmm�m���t��6��m�6�۶��I�[�H� �� H H��e��m& H���{#m��i8   N����$m�t�.� 6�H �n�mI���m�NXHH lz�u��T���Kon��m[�ji2��6Z�Lm�Zl��-@K5��P6�Ԁ  [V�d��[v�  -�����  [E�6ݸ��m��%�$���� [sҒ�l�z�Lk��b�&�FH�k�-�ත��h[�ݓ�
���!�v�� pm��l ���� �N�[�[$���5��(U+�h �X<J�V�^��Sm���[v5�  ��f�������Y>�$�kd� ��|�����a�e�����H2٥�ԆҮr�0�ņM�T�%�n۔kX+:[�n��q��V��\�ـH��ڌv�m��� �91��ڕ�a���vcbP��H3l�Wf �n��+�+q���ְnհH�ڬ�,�5Z��K"[;Bp���lF��z�s�n�]��[*��U�W#� �� H�c�:魶�H 'Z9,�N/j��-���� 3M-[�ݷ 	:m  -76�[v]z�۷:�A���4IM��mݷ���k�m���`�m	 6� � �mi�Z� p j��� pH�v٢�-��IBM�����u�9Y�Y��ܠ�����@Ԁ6݃� m��k�6�` pl�4�6زC�Ho/<�e�@t@�Kcdj�����5�$����ݶ  -����8E6y�n+m�-��WU6nݤ���m����ZK��}o����l��7.��t����8딻l��E� ���Kn�	gP$�N��l-��6F�K���MC�m����{{e�휥-r-6����<��Ht�\eَ6;+5ݶ�\b�HI���[pZ���]�0c8f���ң�-HB��N�`�Y�F� ��$ �vp � ���� ��o�jl֘���-�iY��c�Im �   >u����t�I�o�g,����   l�J��U�G9�C�U��h �@9�knm�m ݳl�-��d�����I"� p6�`��H$p � �u��am�I�� #n�`�K;T�%�8������h��Hhm�  w[&�NͰv��z� ��ͯ`  .���n�n��$6�i�i0M����K. ���}e�6�q6����ݶ[A��l�[i7b@�i%��v�mR�k�XbA��km&�e��[��m[:MJ [@�i ��M��� ݶH6N4�\6�$ �� �d�l�6�Ӄm��m-)n� �m��@-�ր �Yp�'A��[d9�fӦ�lu��L	e�md�BA �I� �m��
���[CZ�m��ۤ�AmɯTzJV�N���l:� ;�����6zݶ[PN�`�1�iy.�  M��e���*��O,����J�  =6ٶ§�v�` ��|��t�-�W�р�= m�زeCb���7:�`l��+.����o���t��.�M�-�k<��(q��+�vN�ؠx�U����m�s�P�U�x8�SAmP�Z�$��E��h-6q��k[d�Xg]3b H      kv��ee�nݳ��N��h $6��XvK(  �mu�m�(��m4�`� ׭�fYD�-�nI+[ۛ[N魫Y�í��8 %�ր     -��L �� ��r�m�  l�l�`�m&� ln�'M�OLm �X�	 )�h�� �m%����)m�� ��t��l m�l����@� ����    �`    m�z�l ��(  m��^�����m�H  ��E�a$�6�O�����  �a��p[@      �hㅴ  �`g[7��w�H6�h	"Z�a��[���� ��.�� �6�;[[l%�GaVu@p �Y@�p[vٲ޺l$   �  m�m   l ݶ��q��  �  9�JH       �	  ���  �kZ@��   �����ۻl����ﾶ�    2^� ��-�l  6ٷlh-i��-�����$     �� :sl  �ל py���  26��$�[p 	��&���nҮ l�۵:�� [[4ؒD���[�t����6ؓ�8֤Ś�R[�@ m� :p��ݻu:������$`ݵ�6H�v�Cs�ׇFŴ��(����u�h���ʹ&�َ.l��Z�v����ȹ�N�W��XHHm�v�f��6��ն�`��f�  6ٵ���m� �e���d    	 ��f� ,�@[N�k6�����  rN�� �v�}�m�K�� �Mcl.كm��۶-�qa������   �m�   m���v��6��V���  ��Im��Zdm� �[�}��]-�Z��6�[dXl��m�-������m�$�`  ;�[]:pVͶ9m�gm�[z�-�ҳi���m��n��  �l����� �l1�b�m��@p[@m�ܑm������v�LV�� M�(�]��jٵ�6���d n�l�c����$n�-��H` ��Wey��Ѿ��h�K�,�fe��8zX��5�vm��L�� $.[$-3m���ߎnGN�2[�� v��YW]�j��j0v�ۖ����۔ؽgQ��i&�4��n�^��:Ŷ�6���mƋ!�m,v��v�M��M�� ����z��[B��N�j�`� ��Ԛ@w�ﭭ�� /SI���v�m  ���` HM���6ؓm&��i h  	 	 �`��\�I��h�lm� �8$$H6�k H M�v�$K(�Izu$t��h�m�ݨ�Un X�W`[c��,��é\�LXl mb�Hs��`mm��t��E�p:D�4I��j��rt�t��lptѶH��۳%'��L(k6n��`�:G6��re�`a��ӭ�m 6��i����h��-�Am  /6�m�� ����u��mm���zY�ln�?�߾�9��8����s+�JI�v�+j�� �%�6�ڶL�UP<� �2ZAڸ	P�y����n�B���m]5�u�-5�-�-�m�"�l���e���6�I�Xj�j����1���m��ӒP �)wM�CE8	e  5�vԭ���� 4TO����' 8�����6�@m�i�	V6  	����۶������m  8  b�J�����`ٖ�J�.��U[HJ�n�I���k�����hʸ�V�  3l��ff�֡	L�5�� �*��،F$ �7����~��-E����U�;Qx�>2 �'ʟ�"�����]A#d@*�{Q"�@`�D ��_��O�+� u�cO��(�8�M���Tk��
b�CI�L@)��� �3�O�E� ш��T����!���Q� �C� �(iT��0?'>tZ|	��R?�=_��P��2� �?(hT"������@
Ǌ)�1�4�Px�O��(T!@��F�@�����"?E?5�8Ch|�@:⪹����'8�M����uC�E��h�8TS��^���Dt���E� x|!�oc�8
\D8�
 ��v��PD��D� Q@�:	W��LS\? 'qN� D��h ގ�	�*�
�D���΄�� �ψ�.9HAQ��P*U� �i^�#)A@M�!��|�Q�,��7��<���H !�����������b�~B�Z��@��kk�?�QUv��A �� J��`�J  �"��($Q��
�bA�X�!����kV�m��F�-��v��ׁ��'@m� �m��5Ty�d�f���R��첵)�+R��$q�+GE�ˋ���,0رob'��ج���;��s+tbp\��ge��^w\R�)�ۮ	��e��\�t\����/���uˮБZ��n$�s��ɗ���;��R��Di�K9�L��K��2��ǯh�|�&��l[F��Oeh�/c#���
'f��5�s-q�K�bݹ� �u��M�{k�����c�I��OKuٷWIrI�Y'E��r���-nm%%��q�^����^"�@�)ՠ��q�^�M�r$3�n���-��aY
���GK(��zm;*i�6�7ZA���l�i�C��*l�e�*N��@���t��٭ �@��5ڀn"�K;6��zv�kiv�`�9�)��ݤ�>�Y�+��s��0b�Emiu�����탶�N�����virY�i5_P��K��ڲ���g8wn\S ����m�{.���tpI Mvz@2�J.GY+.7�]�]��y�vy�ΰ�<�;��75�Ga�jɴt�����t+�qi�vzH�\K=��I��}�x�Z�t�#n���^Kk�	s�U����:n3�����oI�h5�3��@6�RU/6[ �m��x�j���ŞP�����Ў�ngf���]3k�4�඲�k�6�F��n�oJ�MoBmT ����ҼZ�0�bԇ��K��r�.���1���]�dc��e�Ѯ�9K��v���Di���K�'�0�*��c`Ηnk�8CS�������P4��n�6�ZS;<L�i�fn�+��5R��]��{*j���qs��ˬ��d��*4T�Ѣ��-�F��X-8J���3;OOg�p%�V'r��Lj՘5����f�t�A������vUͭ�q��m8�ؗL���b�۪��gv���_�vh�۹n��Ѫ��E�т�h�Kgq��g���?�R'@\v�t�Aw�DF" ��l7��1��m0��z ��G��n��a�^v�O)�e����t^U��Zo��uӷY{U2��l�U�����£	t����nn��yl�WL��������j����l�c�;Bd�=˜>8�g�n���n�-L���WP饶�W`�<l@cf����zVn|q�
U�ϱ�&�`k�a�t]�۔��e��v�s�+kL�:{p�h����m�{����w��o��#�r nx�0<+��y�3��W�`�;l&1ȯ;�1�>�:��x��i`n��0���+H
�MMTQDլ�m���1%Tz���.�zm�h�c��e�R��"�y�h�th}�zD��k@�y��["��$�M�4
���m��=�)�qˆ�k��E�1�m`ۏ@����Қ�\4���J�%�,+,��(J�2�Y�g���j�	�����ɺ2\`��W�F��N(�)1�dX0�g�w�|h�p�9{k�-�s@�A�
���$��4'{�t���7��<�j
�w����X��׶��T�UP�Z*�W�3(�:�n����R]�!�I2a�y�)����1��q��m���$v<��$�F���w�~u}9jĝ69!'3@����m�����w4�q`)��q�x���0���D]�i҂=��;��{<V���\�=sƣ�t��{"�䆁m�����w4oJh���H@�I����I�d�I6��q�oSlp�c�����m����4�0��T� "Љ�!d�DC���T�[u�oZ�ssd�b���hޔ�/;qh������<��l*h �	17����^�z���ҚT(aA��M�H=Ys�ϊmۗ��h����`�X@�)�5�v�ӯmRq�m9�L����'/mz�w4oJh���9�1��4�I�$qǠ^�s~H���>��h���\yLi�V5$�����f��m��Wk�^��Z�iZ�#y�drC@��Šr��ܓ��ݛ�H=LpD��M���U�L�@r;�Yx��`e�j��,g�� ��X^�0�ڜТ;�߿�u�~6�^N�z	���܋�q��6JhN�V�3����t;�Wn)�.�UR����~�,�m��mO�9!W}��.wاȐR%����=�l��jp��X��a��*U4q�����yۋ@��O������Y�Z�6ٗ����$š9��^�ܛZϸ��m��?v��EM��8��;���>�߿~�<��7��)�6z�`(K��%	R�����BۤEG6��J���
b&0�(R��$PH��$г0 )��Q�)��������[;v}/]���%�f^���v�Ґ9i�,AO,�-����W;��`�z�5�m���m�6e^˪w:ø�F��bJ��ɹwF�Ў�a��a����I�����l�M���Ylv��J��g<^s@��[J�J�.7���ݫ�"�:6oE�a�q����m�-�qx�*mR5��i���>���nh�.s�#�gP��D�3uj����D�LM�����Gs��q�.)���i���nVP��M���5��'=����Z݊������~l{M��6z�`z�`�sF
�bf^f~��iU����%�����Қ��ئ8�B��I�X�[��^,�m���S�l��]k5l̗Y235���A"�BB��V��� ���7�ڜg�� ��N�AH�'&6�hޔ�7�ڜg��ׯ���H�O����V��]zk�g�R�y�L�ͶztN7��9��'d�.�=�fv�-�[o��䥠5�w�|���W9_�F��)���!�&5M�&-�m{��3;�p���IJJ�2�b�9�l�7�ڜ�JcOLM��8��=�w4�)�z�ŠU�@�ܙ��W$�0�^V���9J7��nJZ_7z���綦i����3JI���h�.9��sk@o���� �GwW��s�!�0d�i�kAg,M�J8�p8xQ�s����&��`i��
���޻���;�n-��ĤQ!�F3�z�������H�M��䥠5��@Ε���J��E����=o����0�%��jM%������x�h��9-q��)3@�]��
��@����-�s@�;���8E�b�*�� �׋ z�,{M��6M�K�t��`�|�Sit�����^I�f�t;U����}��\ŅWZ���߷� ��X��S�9m� �ե5HWI!��[n������b�"r^������q#�"�JYh⬲��]��׼� s��ׯ ��X�����@��LM��-�������;��ٹ:��@,PYZ��U�<Šz��4�1�4��>}{Z�O��ے���[�����>���2��t��U!qv��7f�t�m�<�a���5�Β��;\�� ��X��S�9�� �׋ �Gh�I�h��R�����oi�9�I(p��I�QG����7�ذ���9J�,vO�����LZ]k�=�)�^�s@�]��T�I�	��	��޻��w49ۋ@��z{rf&�+�$��	��/[��y͵8�n��X �NZjBʩ��b���{9b�ueg��i�\^��t��r���t��=QF9q�ӧK(�7i/U��@f�����p��q�On�cS�����8�,v݇m;�۬�9�v��]�N�h�F��^vs��S��{�u��	��tE�N�лr&�Xv��۩"zֻ��Р.�6�ݕ�i����&��]I�k&ӓ�5�ۉ�^�r���:��U�Ҹ����w�<m&��/nz���'������u���Hy�k��q�U	�AaV6'��x�x�ܦ�w�m����>�Uֽ�빠^�s@��&�� �i�Z]k�=�)�y��Z]J��4�1�6��=�q�)/��K@��^�w�J�ٖ�F7D7!�^�M�v��*�סqu�s@�0x�aH��si�8�(Kվ�poذ�l��r���$cdx
83�7	1J0j�Cv-ϵ��lv��p�c؍i�%�͸�բ�I1y�IUҏRI{�|�<I+��>���ҁ��������?5�s�XS�i�jf�3;������ �1!#Q�PWx&�,x�r���Q�$��n/<I*�Q�I.���&Ю�B'3�J���I%�Kqy�IUҏRI^���Ē�ҽ�a�d�6�F���-��%WJ=I%z�3�J���I%o*�G�G��i�^x�Ut�Ԓ^�-�<�$�K�ԒW����[|������Z$��֓S.k-Cs�u�첣v�sv���d8^0�48.6S��	���F�?I}~���Ē�.�RI^���Ē����]���d��!�ᙣ�����wf���������[o�u��K���}�y�Iu>�<y���$MH�I%z[��H�)5/?vfa�,_�`m����m$8�J�@O���[��-O�c�S��,aE�uk	$HB#!!�����T>�{� �w�����b8~IC�9A����>P� r
��bB22�P���|�B[aʐ-!j�bA� &�!%�l#�o{C����ǽzm�oX�mn��&�LG�RRA��5�Gl!�+��kB5!SK�S��~鉱�^W
pS�5��xp<����|��	T�%D�at;8�l�Ȫ��T:�`�Қ�d����9�m��wvn�oiVj�\1~y!�I��H�)5$�����}ǨԔ�UU]ǲR��$���M�������	�$�[�y�IwK�7m���ޗ��߻�컶��@>|��������68z;�ہ�b0�x읖��x��< �2N��s�)�d��p����Vϵ�J���$�zRjI+���x�^�W��l?,����ԒW����ꪻ�vd3RIG'���$��z��31)?c�.�F�����~�@��~k�����x�]��5$��n/<I*�*Q��c�IcM�jJ���3�J���I[���K�[q�_�Jڨ� "�0�G2�y332�T�:,����Я+�䒑����$��{ߒH}�f���{su$��5f�F���n"b28�v��������[:v�I�a�{"�u�iKfW�.��"N2(5"5$�{:��Ē/JMI%z�3�J���I%iV5b���RI&/<I"��ԒW��<�$�K�ԒW�����͵�豧��"x�q8�5$����<I.�u�J���$�픚�K˓�+b�D�19�x�]��5$��n/<I#�)5$��|�<I/_���&1�8�5$��n/<I)J=�~I%��}���ɨԒ]������?����:݁;���vfh�8Lu�h�+��#Q�lv�V͓��)��1g��
 ���붮��+�=����o[�3�=��&Q��.7C�yM/���w�v>9��v�4�A�fn����7��b�"[�h���9rdI��H�gn;E�[�͌�	8gY��oN��(��Y�[�����{U���i&�,�TU92i�]��h`祸�t�������z>㏹�w��-[u��󄃱v�ְ;~�۷����9�nxM�=�$`w'�Q�m��7/9$�����J��g�$�t��I%z[��J�
��n!%��	�$�[�y�IwK�ԒW����$�l�ԒK����H���x���%�.�RI^������g}>&���w��K�:	ᨁ�$MH�I%�Kqy���w��jI.�~<�$���jI/)V5bŌ$"�I1y�I�I�$������%l�Q�$��n/<I*�DA[0�F�sʼ��:��5���)�n�x��`�Ƴ�q��#�����,o{�x�q8�<I%��ǟ�K�ǨԐ�w��{��q$��ص$�d���QȦ)<I.�w�a�҇�˻o�}�\���׵wm��߷��������?���?>�os���� 7�|����:헓?D%hP�]޷�;
9֒����$��e_	�D	�`���y�I/l�jI.�i�%���ԒK��<�$���9?��$���Z�K��y�Iw;��$��r�<BE�I�$���c��[�;����:ی��X���	��=n�87EĦq���V�BD.�Y�k)�<I+��5$��r�<I#�)5$�[��Ē���xj D�"�R#RI.�,�Ē/K���v�x��K�Ԓ^R�4u�0�	�'�$�zRm������r���B:�
��fy���oK�ԒK޴�x�^�L�j'���RIu�$��w��]m���Kܾ��kRI}��"]Z��]��(�����m�-I%��+�=�ޤ��O�I.���Ē��i�-I���7��$�׎{Z+]�uv���d���W`��Kpd��Q���~|I�u�S3� ����_����$����\��I7�Q�$�u�I�D	���'�$���=������LJzo�ߒJL��RI.����Us��Uݯ��߂ѳ�
�� ��~�߯�{�Q�J�9�r��9!��$�T�^��O��W$����A��<�%������߼Sv�o}�Ms����3v��!Sq Q�D!��Rb�R:��!�*��~�9�m�zK�ݚ�N2(5"5$��i<�$����߇�I+�ߏ<I.�u�K�B�T�#�č�Gc�7n��v�n9o@bzS"YOm�u�ܜc~ǤY��� Hɓ�RK����$�^�y�IwK�ԒK�\�x�^ֈ6	ق�djD�$�^�y��g�d�Rg��IOOV~��_+m^�Uݥ�k8��5�%$Ń��Ē�}�ԒK�Z�ߔ����I'�����;���GLchq�jK�m߯�<�$�?�ORIu�Y��Kެ���F��󞻫G�@�x
��+?~I/���RI{���rz}�I)3ڍI$���?~I'�|b�>XU���.�;l����6JG�y�m��\a�Z)��:[���5n*��w���4��2�cLy��7��;J�XW�YzX�4�r�\+�7�2��9��9xqۦ��:t�vG�|Ӿu�d��]��8ݍ�� �Y7UR�<*�H�8��q&'"g6����K����&B���4��,��.���:���dm�s�YsF�ѢTȨ5��!��1��[cqK����7O']���cuc/�B6ny�;I��q���Z6|��8F��f���$��z�I$��2W�ZK��W�$��[K�6�#�����%����詈P�I���]}���ـyŠ��8Ƞԋ@:�M�l���_���;��hR���#Ɍ$	�&��ՠu�M�_U��%~��h�D<O�%y�p�:���o���x��v����-Q��g�]��n;q#�v����󇇪��n�c�fֶsq�����ύ<�l�s٭��ߖ�u����M�Jh,�v~I�œ�qh[I�����{���A5��Hˆ�ZZ�|/��o�k�p:�C@���[8�:Iuj�*EZ�]]��}ِ�:�����z�۹�������b��-bJ˼4'�a�w�����Ћ��@'Z.U��$Ds �r���@���:���u�M�{*x,��,x�N%�;7<�=7m�K흖�<I�N���>v�-�>���a�Q����XZ�_��)�x��~_vL��!�s��n-�EX�W�YH3+L�Yx���(��RD$�P��}���:�yh[fl�$64aut�V,���� ~w� �k\�P�[,�I%I%
йE}���_���U9)54eٙJ��4'*����9!���М���h*n����YV]�Yx�[e��=�����`�k�Skn���ŝ��k����%����h���ٴ��7
'k1l�x�ڟ�w��Н�lq�.JUUj��~�^�0v��(��h�"�xU�-bH�y�_q�9Iv�Z �h�u��q ��.R�(��m�C@�w�= �i4���]��f�=3Ɓ��`��y����˴�/BWrC4�s4��43����HHb`X�"�h�)���5�!�4��3���;'���XO��c�(�p� ���%S�a��r- �l���Ϸ���M.���D�ms�j��[�2Z�xպ岠c�k[Av�ߞ�k<����+)M�� ~w� �i��m��� ��hu|G�u�V$^e]xh����.�͆hz�h}�l���j�RVReYv�e��$3@?}ךz�˹�4��Z���n T������3B/��-ǐ�?}}kC��NHM������_��@�Қߗ[� ~���9��p��
D%��Θ�q���\1����	�
\	"��!�"D"0�B@�$�B D���DE�HU�@%[
D�҇r��7O5�F?��s��ΟǑ�@�E�d0�CH0`@!tČ�C�jA0N�B	�@�h'������4k��F@� �B!�FE A�jH�$aa2F1��u\�������������-�!@_L��K�
a- �B<R�bH�#,�HĄc#C���>��.�N���r5D��`v�А^�wTc|c
����HY9���TȄ�!&���w�}���oz�o��y`(
��-�� $Uѵ��m�N��` U�­Zl��������ݵ�9f
�����tۜ�س��-�^�F���-�onB���1R��E�ƑoQ�a��]���d�á�����x�㙋�()���p���1R�V*�6�rްnەz�m�1�I(mM��Yz�4�]&�����O�\y�{�zkl��H��Ԧ�v�u��2��L�.R��cm{.����m��W��5�,�l�5bN��n�ve�t�m[-�v����A��#Y�YSB��q[l �\��fy�9� �O���5�Hre{m� ���K���c��ug���9�Nػg�`ݔ֑ewb�&���(ڳ� ��(8�8�v��K ��K(�{c�K�2�Pk�7-���u���}.�Rly8'���(���5�8���'gW6�`6W�'6��u;n��mO��݀.8&ٺWmk��mԨ����]�;If����[�86F�,9@7St���0i��`;k���S`�C[Up��p��N7�3���k�ۍGWam����mNW;	hEjTH�F����24<�r����ZOE	�l ������؛�+��k��v�;n�+U�mu*�Ş��r�� ���o��G�ɂ� �����ڐ���e4�D�P/"�mPng�rͺvA�U��u�Jʇ6�ҭpm�It�Z�n�L����Wf�rmJ�HOm�9v-�c��iד�+mq�&1y�$/X�^ӄ*_6��ƍ�iY��U��F��iWu�K�k[G汘��	V_VL�p�7i��%ړ��0����S�+49�#��ʪ�5���n8� "v;��e.��U+�8x�u��Nv��wd�mb�E�43V� �Ù�VΧ��t�f��v�9�t�F��O�����	��k�vˉ��Zl�X0��N�����Q*��Cfڹ�`�۝M��H\��gK�@��A�K�<m!5�i^T��F`rg���o{����x9��. @8�y����Ӧ '蟕��lE�.�>u1@.pԙ3'�5%���3F��n[��:r�A�zF�����m�)5Dw^� ����k ��e�&�֍��cFx;A��R��7N0�`C��i�ۍ�C�\���i�1u*���n�aȲ��ְn#�M�n���,�v
yU�D��B��p��c�&��)�h��Ü��2�V��M��V�����C�*���vSu�y[&pۿ�����>��m�N�����{���i~�V��V<�J=�M۶������q�'g��p�d/&���q�����hu���hs��)�yփx�dNc$n' �l��Uq#�n-ǐ�?w���V�<XHD�M�hs����s�\���o!�Hd�W+��0x�}�O �R-�gƁ�t��sl����@��|DEԥV�,�T]�~�q���~�n-����;�����xH�;C�e9nlvʖ��+^�we��K����v��cb=���`w��X��Hf���ִ�G)��C���L�bX����M�"X�%�����S��R�%՘fkS[ND�,K�뾻NB��"���IU�Ϊ�CK"n%��{|�ND�,K�{�M�"X�%�{�zkiȟ�,L��,N���f���մ�-�]�"X�%���o�m9ı,O���m9�Ľ��5��Kı>�뷿[�oq�������Άce�Y\��9İ���ߦӑ,KĽ��5��Kı>���K��dO{��iȖ%�b~������tj挚��fjm9ı,K�{�[ND�,KO����9ı,N����r%�bX�w���r%�bX�=;��r�W2��	��q����f�v���w�+F�;v�[���%����N��g<v��mm9ı,O����9ı,N����r%�bX�w���(@C�ı/�������bX�'��73	�2�\52��WiȖ%�bw�ߦӐP,K���ߦӑ,KĽ��5��Kı>���O䀦DȖ'�l��/�,ˆj�356��bX�'�{�iȖ%�b^�ޚ�r%�C��1���2&D��o�iȖ%�bw�ߦӑ,K��?v���P��2f\�5��K��F(�=���5��Kı?{^��ND�,K���6��bX+b}��I���}�w�a�Y)r���35��� �'?~�pI��T���ͧ�X�%��{�m9ı,K�{�[ND�,K��m�Dߗm�q�{��8x�Q���Xk���c+�m]-u�}�7Ϧ=\���ܿ{�"X�%��w~�ND�,K�����Kı/}�Mm9ı,Og}��s{���w���������Q���5��Ȗ%�b{���N@,KĽ��5��Kı/��kiȖ%�bw�ߦӑKı>�|e��5sFMk53Z�r%�bX�������bX�%�}�m9ű,N����r%�bX��ͧ"X�%��ޤ�z���Z��Ys55��K��?�����"X�%���o�m9ı,Ow��ӑ,K���")�D����".�T�1 ł�%E����j���Vk���'$O���魧"X�%���ٹ�K���V�Mf���"X�%��w~�ND�,K�����v�D�,K����kiȖ%�b{;�fӑ,��oq��n�����tn�B뱪�K��ú���9��q��㜦�zd2sp��������.j�5��ND�,K��{6��bX�%�魧"X�%��｛ND�,K���6��bX�'��ܞ��atI�M\�m9ı,K�wƶ��bX�'���m9ı,N����r%�bX���ٴ�Kı?~=�p欔�Iuf��[ND�,K��{6��bX�'}��m9ı,Og}��r%�bX���m9ı,N�]=���G4h��&f�iȖ%�bw�ߦӑ,K��w�ͧ"X�%�{���ӑ,K����ӑ,K��?����d.�ԫ���̅����$'Z�X��bX��3���5��%�bX������Kı;���iȖ%�bA4��;��\��lԗRB��Z���V��I$�sm�Iy���(�{�\��6.7�N���g�X�6��9$m�I�M�����1*U��)k8����Rv��ws��m�زD��y�c���-ӷMٖ�2��i�����o>6a��7mx:�;2t����6ݪ�݀E��g�cY��ʎ�!N<�h�W�y5�'���m�UNݛ����av�v�g7'��g��{�����קʛn:Z�+7j�V��U����kU.�����ܝm�F����&iѫ�2kY�sY��Kı/���kiȖ%�b}�w�iȖ%�bw�ߦ��7�Q,K��fӑ,K����7��P�$�֥5�5�[ND�,K�k��NC�X�L�b{����ND�,K��fӑ,KĽ�|kiȖ<oq�ߟ���/o�3��3������bX��w��Kı;����r%�bX�������Kı>�wٴ�Kı?���3�Yn\պ��ӑ,K��~�iȖ%�b~����ӑ,K��=�fӑ,K�﻿M�"X�%��wy=r0�$̦�k6��bX�'�ｭm9ı,9�����f��Kı?���M�"X�%����fӑ,K��2H{!.B�hөn���ή,<�����q�۶>��-tWl��fÒ0�ɜ=F�،ڪ�{�{�oq�������r%�bX��w��Kı;����r%�bX�������Kı;�t�kY�Mѫif�ֳiȖ%�bw�ߦӐ�_�ʪ㸛�bw9�fӑ,K��~����"X�%��{�ͧ"�������q������,��\u&km9ı,Og}��ND�,K�w�ֶ��bX�'���6��bX�'}��m9ı,N��%�N5�hɫ��5�ND�,�"\ｭm9ı,O����9ı,N����r%�`O��￳iȖ%�bw��y?�L�Ѫh�f��ND�,K�k��ND�,K�{�M�"X�%����fӑ,K$-�~��\!I
HRB~����/��Ms�ӆ�ougl��VUѨ5˓�8-��k�Շ��y�=1�]gC{�[�oq�����iȖ%�bw?wٴ�Kı?~�}��r%�bX�{]��r%�bX�1�=�g���\չm�M�"X�%�~��ki�"$r&D�;�{�Y��Kı;�{��9ı,O���6��bX�'����d���[��W5�q>�bX�'{�k6��bX�'���ӑ,v&���#]<Co"dO���6��bX�%����ӑ,K����Ú�R��3WY�]�"X�!b~����9ı,O���6��bX�'���ͧ"X��*�����v��bX�'�����.j��4[lպ��r%�bX����m9ı,�?{ٴ�Kı>���]�"X�%������Kı?�_㾖^e�5���V��$�:玟X�+I��r��k��"`w�e��<s��l��S����~����{�����ٴ�Kı>�z�9ı,Oߵ�]�Ȗ%�b}���iȖ%�bw��.pѪf����iȖ%�b}�t��r	bX�'���ӑ,K���ߦӑ,K��?{ٴ�ı,O~�&����a���s5.ӑ,K���]��r%�bX����m9�,K���fӑ,K�����r%�bX��}4f�5��52j�ӑ,K�����iȖ%�b}����r%�bX�w]=v��bX �睏�Q8���~�ND�,K�=��3�Ys.jܶ�ӑ,K��=�fӑ,K�����r%�bX�����9ı,O���6��bX�'���C������z�����sЯP��v���ս����9���w9����_�Z�:՝u��O�X�%�����v��bX�'k��ND�,K��~��,K��=�fӑ,K�����Ú�R��2eѫ��Kı;�]��rbX�'���6��bX�'���6��bX�'��O]�"ؖ%���Ǯ\�1�4[K�u���Kı>�w��Kı>�wٴ�K�V"~��]�"X�%�����iȖ%�b~�{��5iLˢ��-�jm9ı,O���m9ı,O����ND�,K���]�"X�%��{�M�"X�%��{�fI8h�3NkT��ͧ"X�%��u��iȖ%�bw�w��Kı>�w��Kı>�wٴ�Kı8��81}ߟͿ81����ہ;��d^�tG:k)���z"J�-ޝl.�e/=,	��jLU�8r����r] �����-�9�i5��t�z�N^*�'����X��j��i�\3�����`4/V;F&�g%����ݺ��r��&˻hIyFk�{"���x�T�D�y�s�?��V��Cs��nΉx��t��s�`c�sFX���=q�:�8N�{���w�?��]�w�m�&�]X-nx�Y�ڮ�z�q����6��gG)�v,1��<r�{�8���ώ��֮a���Kı;���M�"X�%��{�M�"X�%��{�ͯ"X�%��u��iȖ%�b}����je��ɩ���M�"X�%��{�M� ؖ%��~��iȖ%�b}�t��r%�bX��w~�ND�,K�=��3�Ys.�f[sSiȖ%�b}����r%�bX�w]=v��`ؖ'��ߦӑ,K���ߦӑ,K�������H[��k5��r%�bX�w]=v��bX�'��ߦӑ,K���ߦӑ,K�!�?k��ٴ�Kı;����3��XaufL���9ı,O߻�M�"X�%���ߦӑ,KĿ~����Kı>���9ı,O��~��]ѐ�휃pp�D�����/]�\� +V��m����7F[q��cv��jq>�bX�%����"X�%�~��kiȖ%�b}���]�Ȗ%�b~���m9ı,O��=fh�Lˢ�Z5sZ�ӑ,K��?{ٴ�1���]�4��B��@Z$]�dO�X����]�"X�%���ߦӑ,KĿ��kiȣbX�'}�I�$�T�9��.k6��bX�'߻�e�r%�bX��w~�ND��b��2%�}���"X�%��;���ND�,K��7����kD��.f�iȖ%�b~�w��Kı/{�kiȖ%�b}���iȖ%�6'{�g�iȖ%�b}�n��j�-�Rˬ��r%�bX������Kı�｛ND�,K�׳ٴ�Kı?w���r%�bX��B��Nd�f��ԡ�=v�p:�.ɹ�w��=:���rt]cg4�:��{�ۏZv~p
Q������{��7����ͧ"X�%������r%�bX����l?�F�L�bX�����ӑ,K�������!n�.Y�ֳiȖ%�bw��{6��bX�'��~�ND�,K������bX�'���6��ؖ%��ǽs&r�lp��5���m9ı,O���m9ı,K����r%��HmN����fTЮ�|D
���kK5�B\+�	��Ý�:�&��>>@*�0W.>eb/胟�@\ώ��|HSjT�5��+�1I�d��GEMSF �!���YQ�Fl(�GpR��XA �xJ�ù�h���~���'�C")��
D�`Db�@�M�ɲ�G_�\�PC��$�O0>��6.���Go��QS�|,�#�N��EM����!�M��?(������'�~���m9ı,O��g�iȖ%�b{���3Zk�h�ɭfjm9ı,N�^��r%�bX�g{��r%�bX���g�iȖ%�b}���iȖ%�b~3��Y��2f�LԗZ��r%�bX�g{��r%�bX�����r%�bX�w���r%����=�����Kı>@����RY������-�47:M���d�9��
-���Y�|��g�z��n�ts��dIM���Ou�g�"w�����r%�bX���6��bX�'}�z�yı,O����9ı,O{��OkSi�SD��ͧ"X�%���ߦӑ,K�ｿM�"X�%��{�ͧ"X�%����{6��bX�'}��0��fk-�j]\�M�"X�%��{~�ND�,K��}�ND�,K�u��m9ı,N���6��bX�'�?����&L�Z�-����Kı>�wٴ�Kı;�x��r%�bX����m9İ/�A��'}��m9ı,N���z2��V.��kiȖ%�bw����Kı;����r%�bX�����Kı/�ﵴ�Kı=�x����T�����7fT��u�{k����ґ�5����{m%	�=����`���ʗG���Kı;���ӑ,K���]�"X�%�{��[ND�,K�׏]�"X�%��맬�i�a�,�]kFӑ,K���]�"X�%�{��[ND�,K�׏]�"X�%��w�6��bX�'�?x���S&h�]Yu�]�"X�%�{��[ND�,K�׏]�"X�%��w�6��bX�'}�z�9ı,Ow���N5Mi�MY�m9ı,N�^=v��bX�'{�6��bX�'}�z�9ı,K������bX�'��o&{Wi�SS3]�"X�%�����"X�%�� ������O�X�%�����m9ı,N�^=v��bX�'� �&�(f �"�T �D����P-P�5 `�)������o��?\�ɼY�MiN�,kщ� 	Fg3� �w��h�6��/(��c�iV)��X�p�]�$���I���C�k�8#�g��#�JLx��8�!�nl���^�[j�V�ؓ<��.J���n�nEr�T�z�Ķ�ȵU�c؎0��[Yx��:v�;I��9k[���<#��8��śg�"��m�����R���zF�F�2`������{�w{��[�:it�n�c���׆�׵m����7iV��;�u��]w[�T���D�ڝOD�,K�����ӑ,K��{�ͧ"X�%��kǮӑ,K���{�ӑ,K�����{rY�Y��j�9ı,Og{��r��DȖ'}���ND�,K��~�ND�,K�׽v��bX�'�k�}�J[����]�"X�%��kǮӑ,K���ߦӑ,�!�2'����v��bX�'�k��iȖ%�b~�wٖ�-�̒��̺5v��bX�'���6��bX�'}�z�9ı,O���m9ı,N�^=v���S"X���\�ӎa�,�Y���r%�bX������r%�bX�g{��r%�bX���z�9ı,O���m9ı,O�׳�c*�r>�u��Hǳ��m����2n���ےbpc�H^xΖ�x�7d:sU�r%�bX�g{��r%�bX���z�9ı,O���m9ı,N�^��r%�bX�����N5Mi�Mj\�m9ı,N�^=v���5 O�c_8�;w�,No���ND�,K�����r%�bX�g{��r%�bX��x���h���MkiȖ%�b}���iȖ%�bw���ӑ,K��;�fӑ,K��{�ND�,K�ߝ�����i��[}��oq���������H'׽�lI�?w�t��H���{�M�"X�%������ɚ�-���r%�bX�g{��r%�bX���siȖ%�b}���iȖ%�bw���ӑ,K���R���~vH�;Cvc���|�O�
�WM�x�r����t���?N�{)�'Cf��%�b{����ӑ,K���ߦӑ,K���]�"X�%��w�ͧ"X�%��{}m��e�$��34k[ND�,K��~�ND�,K�׽v��bX�'���6��bX�'}���r%�bX��z�֜3,ԆYu���Kı;�{�iȖ%�b}��iȖ:Ey	詭�bg����Kı;�w�iȖ%�b���y]�HIV��Ww9�)!I
D�;�fӑ,K��o�iȖ%�b}�w�iȖ%�bw���ӑ,K���.BpѪkNjkR�iȖ%�bw�7��Kı>���Kı;�{�iȖ%�b}�w�iȖ%�ouߞ�����ى{3گ<�Ը�^y���6�V%ۮL�Ä�ݤ,]���r�jx�Ԛ�2����%�bX�����9ı,N�^��r%�bX�w]���%�bX����m9ı,O��}s5�r[�������Kı;�{�iȖ%�b}�w�iȖ%�bw�7��	�L�bX���]�"X�%��;�L��\&LԹ.f�ӑ,K����ӑ,K��o�iȖbX�w]��r%�bX�����Kı<~��		uIMXfRk5v��bX�'}�~�ND�,K�뾻ND�,K�׽v��bX� ~����羻ND�,K�{}���ܤ��34f�ӑ,K����ӑ,K���]�"X�%��u�]�"X�%��xߦӑ,K�����#g�I.B�X�٣E��]�>8�h8�s�5��l��#�m�NI�J��]Y�Me֮ӑ,K���]�"X�%��u�]�"X�%��xߦ��	�L�bX���]�"X�%���z�Ƶ���4L�њ֮ӑ,K����Ӑ�H�L�b{�����r%�bX���]�"X�%��k޻ND�@ʙ����䓆�S4d�֭�]�"X�%�������Kı>���Kı;�{�iȖ%�b}�w�iȖ%�b{�5��S0�Z��%�5v��bX6'��}v��bX�'}�z�9ı,O����9İ?�U�Os���ND7���{�����������}��ou�bX�����Kİ���o��i�Kı=�����9ı,O����9ı,M�b�`&� "}@^;'�e._Y�t�2d�Z�lh��ʃz�b��r��vN�D+vk��@ӈ�!�ٟ�/���;@{q[lg�fQ��*�w/۴��a�κ\���\coi��v-v�*��Z.�8M�v0=�s����v�
��=�ӎu�(4\��nHȪ��)cncgd����J3s�Ň<NEUv�U�����<[{��C:�!Ws���&���[�Tճ��N�Ej�+?�{�����{�7bN��ݞ��λW^/m�v�1�<�^�9W��!���s~{������	�5.K�����bX�'���]�"X�%��{s�iȖ%�b}�w�iȖ%�bw���ӑ,K�����$%�%5a�I���r%�bX���=v���,S"dK�����Kı=�����Kı>���Fı,Oߏ{,��[��Vd�֦�ӑ,K����ӑ,K���]�"X�%��u�]�"X��2'���?�ӑ,K�����2�N���	����r%�`���{~�ND�,K�뾻ND�,K���ӑ,K�)�?{~��ND�,K���?�kYInh�	�3Z�ND�,K�뾻ND�,K���ӑ,K����ӑ,K�ｿM�"X�%����)}�����K��5���uۮ�x�s]R#�r�ڶq��>Wm��kX�-�^���r�{�r�{!n_�ߓ�g��u���۞�ND�,K�뾻ND�,K���6�"X�%��w�ͧ"X�%���׌.z�I5�5reɫ��Kı>���>E0C�
�O"r%��{|�ND�,K��{6��bX�'}��]� ��bX�=�zh�]fe�R̹���Kı;�o�iȖ%�b}��iȖ%�bw����r%�bX�w]��r%�bX�a���e�	�5.KsSiȖ%�'���6��bX�'}��]�"X�%��u�]�"X�-��{~�ND�,K��oА�E)��e&�WiȖ%�bw����r%�bX"������%�bX������r%�bX�w]��r%�bX�����|�����Z�ۮ�\s�]<9;7��ݰ^�7OWg���n!E�3��k�1�`N�L�����r%�bX�w���r%�bX�����Kı>���Kı;�nz�9ı,N�����i�p�,�k5��ND�,K���6��X�%��w�ͧ"X�%��{s�iȖ%�b}���iȅ�bX����ƳY	nh�	�3Z�ND�,K��}�ND�,K���ӑ,z��b RB2xV�9�=���m9ı,Oo�iȖ%�bx����TѣT�5sW5�ND�,�D���'��r%�bX����M�"X�%��{~�ND�,������r%�bX�݆���?��!�S&S56��bX�'���6��bX�)�{~�ND�,K��}�ND�,K��M�"X�%��jz��^��N��1�9o7�ܙ6�[�&�l��:�q؎vCX�׉�f����U�Dm6��l�'"X�%��k޻ND�,K��}�ND�,K��M�"X�%��{�M�"X�%���|L�Yp�f��s5v��bX�'���6���@"dK�����ӑ,K���o�m9ı,N�^��r%�bX�?{~���)Md3)��ͧ"X�%��{s�iȖ%�b}���iȖ?�EL��=�����Kı?g���ND�,K��{2^[-�K�2fkSWiȖ%�b}���iȖ%�bw���ӑ,K��;�fӑ,Kz1�Ah�$ �����@剜��˴�Kı>�{5�Ӣ�,�k5��ND�,K�׽v��bX��?k��ͧ�,K�������r%�bX�w���r%�bX�������a�]K5�5�C��D�v��k
�9��k��s,�˚�$�t�B��2MY��]�"X�%��w�ͧ"X�%��{s�iȖ%�b}���h�bX�'}�z�9ı,O����4j��&�Mf�ӑ,K�ｹ��ı,O���m9ı,N�^��r%�bX�w]��r'�S"X�݆�����CZ&�L�5v��bX�'�{�iȖ%�bw���ӑ,Vı>���Kı;�x��r%�bX�=��Y532S5rff�ӑ,K?�D�����ӑ,K���{��9ı,N�۞�ND�,��~�ND7���{�o7~;?���0@�����X�%��u�]�"X�%��kǮӑ,K���ߦӑ,K���]�"X�%��j�CP�Ĉ �A
� sH�����'�ؑ"�BmZ@d҄��]>a	���\��5�߶=:BE�ȸ�2�:�D~SHH��E�� %JTp޶�K�N���+�N"m"@�"ET�`HE	6*���(��"�Fr��H EVVD� ������(�E�_�0dS|��	 A )-Dʤ�2�ȝꌐcCp�)���GR/��!wb��/1Ȅ �_�1 ��F	��*h�"E`H����aN�>�_��R|����i��	��6��� �-�����\tj�+V��=n�@Gت��V�b*Öɫq-��A0]�*Q� �Q���)ݬ�{870�ڷN���%�\e��ۜV��W=h]	�6���;���Vls&T�Ҷ���]�L���l�z��v�ۓ��
3�K�Kf���H���Y�:�M�����7r�94��(v�����]�l�N�����9*���E#E�l���f�pK<�zCK�l�����f�efU�(�Vc�<����n��8�r��ݺ��tlT�M�ڞ�g�ҶX</n�$��nXW�lؗ�#'q��Ͷ{S��ء��!Ց�荀�6��0����'n�*�����{8��4��9�[,f8y��p�nIl��.���:�m�.m4.���]>==v�uMby�'2�Ë��`L��n3u��J�I�u:�ƣ��[J�	�������nWb�[K���m��gd܌\-�Ѷ��[Z�U;\&�zj��Qͅ$���sٝ�H�f�Q�����An�peݘ��N������ju��k��KÎ��m�.��y\��wY,�9���w'�:��TC���0 �j���9�^����lm���`L�.����*���H]R�\�U��gn6� ���oMvɵ�+��b�mD�kʀ�U� ������6H-�n�N[m�&NT�	�\&I�k$JԫHO'�Q�;ZK��Ρf�@�㵚ͻq�Bv�٫���pvK|�&�w4�5���`Lg3k�'FF��!���[@ۤ+V���Pt�P�g�WUi�]ȾW�b�<<��Lk��n���{\��M%��Ei�ۑ���<�[�qY�k�|�=����i$:�X�G8ٶ$ڶGA�ܴ
/7�٨�.ZxZ�zQ�[:�&�*�Nw����P �ل]���L՛��|"��k]�s��]��u�`W���3��|���ꄙV�p���; ��wm�]K���h���������u��t b�*1���+���8)�a�'���/r�n�`M�q%l̑g���セa^Ʉ�J;ɪ�rb35iwk �֫��5�.w6��"�gm�㞞ܭ��m��N���c�^R{�Ŏ���5j-۳6R�;U�����=�ӟG[�.�Aݓ�rǁ�j��R��ٹۧh{hѵq	��t���Je]Q��͞������!kN�uwV��
ëtF�˧]�u�E��3Ve�B(��������YN�u���Ҏ��ݗh�nq[��\[>v���p�ר�ݷb�&�v���~oq���?~׏]�"X�%��{�M�"X�%��k޻�DȖ%������r%�bX��?����e�YufL�jj�9ı,O���m9ı,N�^��r%�bX�w]��r%�bX���z�9��"X���f��t]VMf�SiȖ%�b{�_��iȖ%�b}�w�iȖ%�bw����Kı>�w��Kı?{]��f����dշ5��ND�,K��~�NC�9"X�����v��bX�'�{�iȖ%�bw��������$/*���e�E�j��&���Kı;�x��r%�bX�w���r%�bX�����Kı>�w��Kı?�?���ZS����4m�s��^D�:��_*ɮz��Y;s��b�ۓ�Y�\�����Y��~�߽�7���'�{�iȖ%�bw���ӑ,K���ߦ��D�DȖ%����iȖ{��7��������:��r������%�bw���Ӑ���X��´#Z0^�䪪D�K���6��bX�'�׏]�"X�%��{�M��{����w��������g����iȖ%�b~���6��bX�'}��ND�,K��~�ND�,K�׽v��bX�'�{~���J]L)�Iu���K�䁑=�����9ı,O����ӑ,K���]�"X���{�M�"X�%���}2�K-�˫2ff�]�"X�%��{�M�"X�%�=���i�Kı>�w��Kı=�x��r%�bX���K��{]Wl�ҥ�u��N��K�g�Y�h,<R;�ˬݴ��tg{uU�F�w��#���"�>o!�7n��r� �����:���1���MG��t���%ʋ@����ݶ�K��F*��0�T\�7f �4� ��
P4H��"�D	R�
���������0�Y.5#x0�1��hwJh�V��t��k�V�r��1��8���4�{�����E�~�q���a��xk�c"xb	�����q�t���Ɲ��i���;n����y]D�[�gx{6x\sw�@���4��Z��+�	.E�N̅b���Wj��hۦ�r�#���"�?w���URC�8ZZ!+\"˻�Š|�C@n�ZNUs��]�L�{����;��;̼�VZ˫\2�0��9T����y�tօ�>����@? �Q�D￵��6�ί�NLX�0aQŠy�)�V�s�svـ7M��B��վ�%~EI{i���]*��g����s��d)�W��n6{�L�9ɺ�?�����t�����JO����Ӏsvـ7M���f�������P]��*�\�ݶg�Q$�r����Z}IvL�vL��M�\yWsT�U\�UV`�s�svه�	BJWdˋ@�ۋ@��8�˥v]�us�svـu��86����/�ߍ��|`aB�X)ޱՀsk\�ݳ �� ��l$���~t���]Hjٙ,�̎kY�Ü����鶍қ��O8v0����u��r.u��:�c���u��":Y�7va��l�eײ7��u����X�p;K�h�½���#��V5�[c��/$��3�C͊t(�n����n�s1����4��q��֬���NĎn��9+Aę�sem�Tk'�$ �-=�9�z;,"���Wl�S�FY�;��P\)�IyL浬�kmm�ba�[��r�v��rZ��#�2�ZH˻F�Ŋ(!&�
!�H��/;��9�f��g�(�""!.�?}u���>_�G?H҃XF�Z[)�߳��ďm�\ˋ@���[�W+�Ď�j��Uc�cȆ�4m��c�O~K�t�kv�T�jRST����򈈉�]uhu�[)�y��/r�q��P]��EU\���0(����ǀ{�O�ޱՠ^V1�dx�3xc;.S���f-���RVC=������a6ȜM�L�I�hl���S@?BI/��]�o��l�'�W�$�Jf�շ57$���f�"Ъ�5D�s�s�l�5�f}$�U~��F�(������/���-�zSG�u����M��*h���($�$x�=^�U[s����x�?|��嵠�,���55��C@��hr��͇�;&\Z�w�y�R I�އ'��/��קF5����mrOD	��c��E��n��x�V����m��~d4����>���s��92���]�B��*���;���|�)�w��B�~���rCw��9	/�UC����)6ax&��-��Ɓ�ڴ���B�V(P�.��'�ـn��`���X�⻫��1+�4%s�̑h��hu�f���ٰ�>]8�-
���i]��>��4W8䭇�;ِ�:�ՠz���,�4OɄR?�q��h`����eXmՋ\^��eʘ�E��N���m�lO�Uv�f�rVC@���:��������P�	Z�J˼��@����p���RC�"�;ِ�:�c6s��]��,�f^r������h��-�l���䦁��M��*HX��I^f-�J����쬆���;7'W�&�
��@���ܓ���]�Eh.U�ـkjـ}䫕�O�>z��w��4O��j�b��+�Hdr����׎$;u7���+�nz�=�}m
��:�\��&��6�m���&`��7�l�(�\�~�O�o�q7���p�:�V�������� ��f|�%�B�
��dOȯ�I����bWx��x�:�i�q/��h\�@<e ,�Yt�Wha���W�H���hv���9��}����%��Bm`(�c�(�/Jh��UUr�=����yh��ր랪���;v�w�������cnϥ�[��"e��Ԏ���+{>8p��Zר��l,e[nS� �2nv�VL��Gr�k==&q�s�ݷCs��2t��7�
��7N�6��6)í�83�s�.�ip�H��6�ء�.�6�:�T˭/�+�	�W:&�77�&�w��:'������cv��pa�Xs<M�Oi.�n�ٱ��'t3ϭӛtm�����������QZ>��>�	L�k-.MD��^Ag;::H�ٮ�}r���|�He:$Jf�8��Wvtmo� �ֹ�7]˟�""�=�ύ�e>C�8�1ē�-�_Z�$71E�}C@�����s���.�}�I�I�E!�[�_-���ܮU9�/�>����鎮��A�F+��[>�!�9r-�w���W8����BaVEx����.���h�Jh�*�/Jh����<�����v��f�o0�l�5��3�C��e�=2pį��������ݟ����Q&���|h�*�/Jh]�@��L Q���
C@�U����_�����A���(~�	DJ�ï�K��?gMˑh����U$}Jj�+��`��3-��]���r��}s�@��Z��;s�Q5�rC@�M���f��\�}�߽ό�?��',��`�C�-��M�""M�'��;�~0t����.�6�t�/k�8��K۔�\�Dv_PS9gg�LzۭZV����wwu����η��x�� ��Z��4�ՠw�w4o���I�M���@�������.E�>���~@����
�+�v�h�ʪ� �v�{�Ԛ�� v�h X�)�;J�f�I�M~b�	"5iF9���5�@���3dc (E	� ��*��`����bcʡ��ʴ��{�I��	��]��(���{R$�$�bp@�Bi#���1�$b�C�$�&����a>�ic'��N�ئ@!h�>B�Ұ���S�N&��|�������DQv���'4;
=����IS�˞N��%tR�L�WV��+2�+Bs��.9�@󘼴ץ4���`�hō�N,�n\�B��F��|t��׀su��=�Jb?\�$��#A�&H8p�zi4�:w�ܓ��N��ܻ͜<�/��(\܀q���S4U��� �w� }o�׋���b�hZ��8���k䆁}�~B�����w>�����BS&��>�,��`�Nf��~��/�X:��x������V�l�%�sV�=
�k����_���X	(�DE!ۇ�l����7$��\x�1��0��Qhu��/���;��`�N��>J������F�\�엯��c��"��l6EɴS�㱺G��;7���{��?nw˱8u���{���׋ �ju��v��N��Jj��ɲ�`�x��""�ݩr���h�ok}T�Nɔ ��,J�UL�լ�R�X5�0�D$�{��f�����{�%*�M���I�������g���b�;��`z>I(P�^L���~̻�^X�Z�/3�m�����k��� �f�hJ�{�<���� )�~LRb�&D̸�6"s�i1l��Snܕ��3�9ӴUӘ��gn#�㧮;68����n��ɷL鷛��wF���;/	�B�����&׭��u�ŒQ`��j�Sg��3ll�әUw.դ;&=(wa�����b�ɹ�nyݐ�m��^�su�<5����f��9ѵ/8�\�meb�"Ʌ���]e����!������Z�؊��{��w�0|��nz8�	Lmh�mv@�!v���4tF��������'�w��o�Mr��3^��x��!�}�Mށ�^3�_�v\�@�\��2cP���8h�V�	�����,����ܓ�}�M�U_�En�<g���
�U�F+�Z̽�g��m��sa��R^�_S&�d�Ib�k.�s��9�����:���>�^��YM����:<M��R8��;���=
!B�s�W ���u�s�Z��3x'���ch�0c�O6��R4�"vSy��۝oo96�l�z�����b�<si&�h�V�޲��ڿ���:�6� �E�Z�Ŗ��v�/@�����2 ܕ���;�����������@-��$��&6WV`nـw[Ň��3��ެo��@�_\�1ưJ,���n��R�`nف�
{���-yz.ժ�.&�&��������� �����n��5q,TNĤ���o"��#Y:^ܗ�mm��g�Z۬��v5�cېsѩ�'��2	�jG�{l����h�{^��? �����
���,B��p�<�������G�h�)��Ď�1�\.��E�Xe�V�ܛZ:V���Ja	J��l�;����f )�,m	��~��E~z}�����=UI�?V��]%��+K�ĕ�,������~��7&ց��Z� �P�5��*�I6P�≪UW3�v�ʘ���!��]Rhiu��	w&m:6�^�=ϣ��I#�㉏q��:�nh��hz�W�Z���}��6�x%�h��l�Gݴ��[�@��{[�VbG��}�~�&5	�B	�������Z�ܤ��Z�mh}Վ��輓 ��jG�Z���e4z�hU�Yf���B]2��j�_�P��-�s�>��<��zj�f�V]��Z���ʑ����N^�����?�?�\��&����j1��,Ν砼�qs����8�o#�^#�o9vl𠖭+��9��}�]w�7}jUW��Xw�������`��A��Л��{�u���Z��}{Z���]�J.��m��|��@�|@;����k�z�U�܏�4Ӌ@����ok@����	�M�@i�EŏQ���!�ym��=��Zs�8�`��(ZDwA��N�l	ܧM��^i:)պP.�����	-ޝ/]Q[W��je�]5khE�Ue�L���3��s����0����D��m͋nz�v��'�ku�L#�]�����zs�psH ��8k�i��&͎�un̍�����nN"<��DKʅ��������;q��yM��������eh����� �ծ�Y��&�ڍk5t����Bz"r�w���{���Z;]�v��1cO9j����;��v��i����l����-�x���ܓp��dơ?(F��@������h[)�ym��;�K����2$Ї"�;�U�yl���s@���o�^����	�]yZ/ux��f-��x�?6���q.��Zv��>Uһal�WV��X��*�ꪫ��@p�����h[)�^�1b�ō����{����h[)�ym��.vT*ŲF�PF����cO�֞\iM�.��]vb�j����K��n��w��v/�e7�hL�n/ �ߖ�岚����U��[�I27<Hn=�e3���F/(IV��,����6w]`�(G#om�h[w4x�����Ěn^����&���u4�Me�ѿ �TC�3����ܓ�￞�岚����V�O��ƪ�(���6w]`(��Q��������}��ց�=Q],ŅٗA��뛣n|:�0�]q�%']n�,D����Ӎ.��<��D�8���=���ym��=��Z.��W���	�L�bW�������W*���8\��"�נyl����	Lx��ci��h��v�I�������JCH*�IH��N;�gM���P���5}
!%��/���ŀot���?�21��]��[)�ym��/RS@=:���8�x�!�� ۶`B�IG�BIB߾���}��h���'��U�2L1��m��'A���F5�jM�6��A�R;e�Y,��3��������6�<��s@�IM��w*���U~A$�hR��Xeeqa����c7�z�Ʊ��$��okg+�����WV�X*�2�/����f��s���_I6���=�8�T�PM��r=�)�y[ŀ=e��
���BIL	&H���_"	��}�nI����L�Y^4�&$�ym��/RS@��^�m�������\'��(������o�G?Wiv���b�����^t�ǋŶe�u�b�J�Ю�2O���3��r���mh�b�
�ᖅV^a�hʩq���!�7׵�>���r��2K.�Z�^f]ҫE�^�$�h���/RS@��z��BH�"F�Yj��W9�#��@���z���U����@�/ORˬ��b�,0Wx���`^��v��x����?�C��??=��y��s F���>��Il-e���SJC!�*}ϐБ1�Ii�#!𸹎hТ�F(4��Z@	����t�'5�&�t�����0� }ut���DڃCD�p�x�5�-֤����� d r�w{����dYh�lm�n� 6�am-�8lޡm�`8��lz.�1�8�L�����v�B���"[��p�#8R8�-�T9:�J� �Q�{vj�K��ʼ�[���nҳ��# v�I-��IG����VĚ;봶y�;��r[���)tK]�kl9(���&x�3J#kj�[[f���ְ���V�v��.TIE�N3����EN��GD��wċ;T���N)"(���de�m���9�'[5�*�$$6 8��g��]��d��1Ԙ�i	��c<kfX��8�{e⶞ F퍮T�5����];۶7H��a�Y2���n����'�[.�WOlZ3V�A�G��x%���p���#�y��]Y @3��+J���u�A�6㋉۞YHe�l��4o;f��q�LG��{sӄ�T�k�olѝ�x��+H��ջO��x+Vۮ�q5�Ҁ��Ց�n�].�b�s�,�S� e�\�A�Z��0�;tx��H焀'l=9雭��wZ�$v�ycq#���v{;!k��yl� ˘�&n��<q�e
fͼ`r"�k�)��7Q�:Yn�8Wm� f�$�V���&x��.09К�E賌��j�d^�͋���) ��WWE���Yb��SU�%&�^Zڪ�,��RK�%��6���Ń�Ku��R$6�[eܹ ����J�OLI�����Ib�U�	C�
�m�|Gt3��#�m��hv�.��]�\ۉ��v��4[�a����U�6VH֫�6��^cMJ���8�dJ%^��/	Ʊ�^:��*�Eݍ�:��]^�*�1�G�e.�q���`f����v΃�6i<�I�>|Fja��y�̛N�cM�-��k���$m[�,��j`�cEq��g7=�*t��m:g�`�pcR�Hہyڃdb�ru���ݬ#q-RXx�\�n�t6�m]������rN�a9�0u��S1dt�m\8k�٫�,W:_S��]K��ǂ�?p���A������7Q~v(�B�"�k$D� �>t&!¨+ۙ��q�s<f0Ə��r$s׫rӗ�a+Ӗ18Q]��$��k�n8��c���m�6Ύ����6���ƞd��ޗ�K��e۳J�0ю7�X݆��vy��=��q�`�w��t����s9�[�i��f���YɯVdu�]�cq�kw/6fs�;M�[l!&����
4h����J=;�wb�nl�r힥^���Ȧ��H�e�e������t��y*hѺ;vKF�;9nk�zz�Q���ipR9�9��U7��]i�u�O$;��"�� ��u�7M� ޼_B��DW��3Ɓx˫�+X����^��78z�`Yl��u�����]*XZ��һ0V+�Z�mh��h^�@�ڴ���0J0y��V����qG��r���ʪ���رB�is��/0�4�]��I�/�H�ր��f�9NW�;�ߗnù-�QMPj��y�ܽ��g�/ts�.����9��w���[��֧q2�J������Ӏ7� ��ϒ��!�����O�G"H�(�rE�[�VqB�P�!qDZ]F��g ��]`�k}�H��d�.����8��]�hL>ZW��-v�޻���^65<X�M���@��z�ՠ[�sBr�sTZ�C.�+�XZ��,����ց��r��G>����@i���<?����q��cj�q:�6�M<i���]���)�v����ԏ��������,Wx�ޞ��^&��]��V���܆	F#�Bnf��,��U���ՠ[�s~H��/���V
����@�9z��W9HA�
I p���K���$MD� D� h)(���d"�>���f h�t]����R�J����_!(����8�mh�f��Uz������/V^fX2F�DҐ�-빠[e4
�W�[e4܈�A��`�$K11���6(5��:�����y^�d-�+.H^���u=&�� ���}���*�^�m��s��H�ց#2��Z�y�.��4�]��$I2�mh�f������-`��3̽I�����ܮs���!�E��v�%t�$Cp�-빠[e4
���y��F(�IZ����v����)]!UH���[e4
�W�[e4z�h��q�]���b�M��-Բv2vcv����vۧ�z�����{�En�ma-�C��s����G/@m�4������I��*�_c���D�d�7�m��:�ŀ6���Y��B�*���W�]�^Z���4	���M���Us�ʤ��^�$�h�}x,2��YVbĮ�'�a�5��mhJ��.z{����x�?��r&�'���W*����sk@m�4U\9(% ��,����'�Ժfe��Y�4�۬���"/\䱋^^�E��-�]���d�b��>4d>�/g8�����&�N�\I��cq���m�.����v.q&ٸٝ:�yp�\�ۡ���a�w:eG˺�q��Jm:�Ƹ���uGT�]��d�&m�������J��qu�2<u�%����N,�n���;�=H���[9/[v�s'<ԗJ�Vv�펧������{���w�cv��1]�,6f�lx�)���k=��\��\��9`.<u%�"q�$8���>����׮�m��r� j9zʺT��)+�v`�Wx��w4l����z�ՠy�LP�፡73@�e4
�W�PQ܋@�ͭ��j�is�^fa�4����ȴ	���l4
�_b���5�Ǡ^v��x��ـ9z� �.�d�R��%�ێ��ٻ�km�����n�XT���ݑ�]��Y��Ļ�GN�l�M�I��������h��4�����;�hB�ĳԫ��E͓Uk z홉A	L$�%I,L�uz��Z�w4x��
��wB�4�]�������.��������h�QF����)#�/;V�o]����*�^���2�,t+���+�-���W9\����>__��yڴ(v*4�Š�7����W���E3!1��p�׫�:���vދv�s����a�F4G�6������*�^�yڴz�h�"U��y����뽜���RDw"�$sk@}e4U\U���$o�&��/;g o^,1d*H�)I!%�\�]���[
z�lBQW��� �:�7��fX^Z��^-Ur��R��ՠG3�@��z�j�<��"x�!s4�S@��z�j�-빡���O��&
�q�AG\u����׶mme��y�:']��Ɓ��q��{���v��<�>9�"L��|��=�h���/YM��(�W�MBA��ιƽ�DU�Z�<�~0�ڿ�%2q~�pO�&&��?��4�S@����hz�2�Ǌ<14UU�$��	*��s� �_���78N�򿔦'z�w�䟾�,�i.[�&$1�!�U�W�^v���s@z��B��kA>�U�MґU�Uɫk�wS)Z;I&M���I̙�m�ͧE՛��ww��>��sR��a���������g�^ր����.�z��0���6�PJ8��]����*���/;V�g��ď~������<�Pm��>�O��z��h޻��G��U�~�@N^�z�j�/���'9\�Q͆���Z	x�	Z�0�=�h޻��)�U�W�{�w����� n�`M�vm<b��9Ćm���]�]�{u�:�nݬ�fci$ҫ��h�֬���A� sٽ�=ȓ�sK�m�W.��pjge���b�Zw.�Ӂ-���e���n��)�Q�ط�8^�X1�g˼��pK=�������Ͳhٷ��?�m��VCc@Џ.6y{I�$��h���7nl��p�l����7^�BA���;/2m[��8����K��[�&MS52\2d��!�B�K��W�Û���S������^N�*�&������,�`^��DDqw"�>�ʅ �
�]����`u���s�=o~BJL��b�
��+,���@��z��(��QU������� {�]U���E�Ǡ^v�����)�Uֽ��'q������@��,��I}���O��������������6x{��]�</��l5� d�n6o<l����	x�:;+p�8�E��h���*�^�yڴ��h�'�U�`9x'��￼�xT�O��E@�_�����'�ͭ��7��URCd]+&
���b�#����֒��s!�9r]�9_ӹ��2�s&��s5w'��2{���{��@n�Zv��?u�2�Q$(���$�h�M�Қ���w���W*S��R��we,.i8��oYy狷�Ʃq����ǟSͰ�F�O���wd�=_��~��nHz_��h�V��w4�S@=��[��<�G�<�Uf ��0�^,�`�k��B����?�D�H�iA%!�{���[�a)�櫄�l�hHG-��>eO�	 �#�V��KVh@��f����,�-Cx}Ɯ�-pB��Y��NM�$�0�-��8�o|����� Xl�lv�P��D����;˥�%�1���4�� ���|o�����;�C���0x�3vXXDa�Х�)��]�������ee>�Dy��@�+�w�� ��a��?�? �G�E��^c������Z��7ԑ%�R�V]X�YI]���� �k\�ݳ�Q=��,�6?���E��篪�:�M��{Z[�h�HMJZY��.��帝qF���S
�J]n�h�x�8��N �iwlayz���Q~������}��u��5�g�>Iv�]{��6a��%|�x� �����w4�S@���h���/�e0B�MbNf��<f����4�K�d4�����;W���\�bE��0��\�)}װ�:�CI9���ܞ~��E�� �D��ki�}E�$Mc�Xc�ㆁ�YM>��F�}�������f k&T����}mW�oI�/N$�mѷI[�Dv�I�=��#���hŮ�6���I������_v��YM�zS@����n��őՊ�Ŕ��hu�6W)#���h{�s�#�H�<5��<��'�����;���c&���`�Z�Y�����M͆��\��=�S@���h/O�ز�O�`��;��$�y�<p�?N ��2I��~P�ĩ��4L-Y6n�4*Y�C-����H[�̹�>��a�^.��3Ҙx��p�a�9Ry_��cy�[M��mOi���q�U[�r��n)88YC��.�+��v�"X�ɵ���,�x���U�R�mn�n2+�5K��2&�ҡu����\`Mf�&h4nm�:��[j�ҙ2��.�@�E��xlO$�9�%�n��p����J�h�$,3�s���ni)瞖��: �?��'�.�l��>���Enݛ������};/^�+�t�/c�d��t��ې�قzݶ,�ܧw��������9��8[�}���,|�5��/�1!���zS@��M�z�h��hwQI"k8���q�@��f��Ň�BJe�{�w� �]�dq�F�D1)�z�h��h{Қ��h���cY1d"�;� �o�Q���o�~0�d�����)���4��C�I�u�R�Ϫ�:��vv��s��d8��n�`.���̜;�e͕5f�v���0�l%�$�����>�]]���R���/��]�ҘD�E�A�N���B�
"�(J����`��Xv�������.4�6A<���YM��X}
�3����7޿��"�R]v���BW���r�����g��e4z�h�S��&�蘐�䆁�ڴm��:�M��h�$^7n����s�5v�eVw/k�����9�g�vvݹ���a;��x���Ny�쩩������5� ޻g�%
$/�����ra��&�b�-�Fl�Us��!�9n-�}kg��Uvw�\�$Z�Ub�1bW�h�<hw��ʊ<�"'�AJAA_��"F&W�\�p|�� }��M*u*kr$Ĝ4���=���:�����M�QG����$N-���UW{�>̆��}k@�UU.ƻ=������ٮ,���i��4�*�r��t������GkR&浽r<.��ȼ�gƁ��M��k�=v��]"��!UL�]���3�BQTO\���yh}�o�#�!z����+��/������:���ץ4u�6�)��5"��?g���СW��}8���0{l��	��H����X�$��
�<!f� Qc����rO��_c�L24��)"�:�M��_��x����:��@��"0���d�&�����ez�G,��w�����8���'��%�J��~�kw@J��r~��@��ZW�hl����'�U�ȓp�:�V��}V���h��<�#x�XX��E"�=���:�3OW9�s�˹�4	�����t�O\k'�'�ȴ�S@�Қ[mhz�����̨QX����I^a�u��{�s$_��9z[�h~^�2 wN��䦤�	���Ùq�1�
nѻj�����v:'��b�[��Ų�2#k�ۋ(ukY�Y�ؕx�l������A�hƳ���)!ո��.aؠq�C^DN������3��͞lhK^�0oRջ�Z��E؆��܅ct�q]X��|�w6ٛ�5���.��m��%���,��a1����x�u]��v�k�Xo&M�-u�����Z31�ݸo��$��3V�5�I���<������v��}]�v9�k���;�"�>�f9�h�]�+/30`=s�����8��_�H�ɸ,�K*�fZ�t�^-��{9��]�{�Z�3Ɓ����+�I1d$i%�@�s@��4k�h^�@��;p��<� '3@��4k�h^�B}�߾�4��l��p���I�p�=�ՠUz����ޔ�=�R���خӊ�t������X���L�OnC�d������Ҹ���	T1���>��;������_�v\�@�3��J��.�����gW�Z�����\ύ�r-��{䏻2�Ee�Wf*)ZB��vd4����)(���[�ۚ��ՙG��m��ػ�qh7/@���h}8\s��M�d�L`�k�ԋ@�����s@��f�Z� ���0��ʚ)
�ʴ�v{q�!�[�G��L�Q� 3v��f�y�wfdOV�@!#ň�9�}��4��h;�_����z�%2���Tǐ$�hِ9��@��W�w��o���#��+����J�^e��rN���n~�X�?D�"$� ��#VH������Пk�훒~���܇R��,�k&��H�*����X�`}���)���p�G�D�4�Q(������h��hwW�{C�Q��4�b�`95��ɣ)	���`��3���ϝ��|����z!�v�|�	�'3@��M������������̍�26��ܐ�=���W=��r��)=z~�ր�x��$5o��bx��h+~z{n�}����Z�خH��<H��̽s�\�O�~�vd4������$A'�� F���9���g���Kb�<� '3@��M����������슥�#q4%&'Y�3%�S��u;^�m���n�=��n�pt/�(�1<0x9bN��Z]�X��^�
䇵ߌ��uTJ���N2H�Z^�z{n�_z��������*4�Q(�q��{Z ���%W*��e�����|�F�l����������mz����kՙ�dm	0rI�w>�@��z��� ���.<�0}�bHF�A���.���Ebƭ"R�TG�s�.����WB�E�PN�@Nb��1UѬ� �*H1L ���8�$x�o3�8p@�JE�1�(�#�@)��}�u����pF`�?1SNu��3\�ky��a�ϭz���<:|����@��� ��YB���)�(�b�����{��׽ߩ�t}���$-��6ٶ�	-��-��m�m�	�-� 8��c2f
�mzMƎ��؀@W�z�)�X�cf�v	�v�Bf�3;h�,�g��,fj�xL"lu�G"��2���Y��\�]�i9I۳uKz�N�M[",�Uմ;v��I����J[U��q��G����ʏ���g`�Ȁ�N�ڔ݃i6t��^����B7:�:M���^����˔l�V4?8�Kv E�oF��6���M7��(B�.m&�gQ�ڮ	n
u��mƎUJ����]5�׭�H]�Xm���� ��DY6�����-�euX#�:�1B�mF=:m])��v��(����\��۞(��c-;f{k�+� �`���w6@;���v�F�e�^!^#,n҆��ܐ�=[rWPd	�`:�n���C8�P<�9�k�t��
�k'&�X�v�:��N�Y6m�^�����J�ۯ.�nZ����V��z[��)c:��6�m���m�rҬnr;;���v��]���'n�wl�`�td��@\=��|��/ �	eq<ݲD^'�GA�I7}�����5�׉4˺�J�z��z��m�3dΎ����t������� ܗ��S2�M�5N����A�Xk9v��m-=�؝
�ck��۬@�܁\�t�ip���ZMͻmWB[)%rַ�-�D�Emq�m���R�ւ�֘����iֶm�c�(�m��� ���K��p-�q.�m[[�n/J�Rm��Rqg {6��c�/j6��pu���Y�6��묎l,��i���"Yv�%mK8�kd���d6�m��n�jd�m�Ye�T�rgNc�G�P�,֎�lݓ<g�d֞�ܺQ��7�5Xь096甼d1��
�77m)���e���-I�q�P����mr�@�T�Qx�jy�h쳏h�:�`�k;;]��lK̕1R�i{=.�e�8t� ��9 �HN�s��m��M���n�=�}�~�^�h���f�	݆��k��v�SJս�SF�n�in��D�)�P����v)�TD�=�PR&�n�
�Q���4�@!�8���D�=ڈ4�F�-���[���,6[��[=lM�[]zd�rNS��B�)�z�Y�D/mf���۹mb�:�N9�Q�9��o���~x��8y�����;��u��l��n1��p��n�۪��L$���!]t��w��k���E�ˣ��D��ۛ݉�T#S�u�v84:ySg9�qΎ� ���zex)�q����;vsi���;Y�Y�sP��a�%�����"��o�K������g�e��k�ʙ/�ۋ��]�0�P5�X�n�6����{�gшM&&�bjE�������s@-�4��h��8�d�28�z�����h�����{��W��vz�bUj�B�@]����}��� ݭs��%�|���}$���7)]^Z�ay�`+�@�o�h>��?6��=UJG��%>#lY�i �d�H�
�W�f{����<��r� n�Z�l�J�,�g����s���d捊�Ws�/-�.��m$[����>�nWȈ�,�����߻@��M��Z]��ה��ɩ���%��w��v�/���f����oSz���I�����9��f��@����՘�?i$�䆁k�-���-����h^�r�ҵ��')Kn^���k@<f���Z�=��`�`"F�Yr=�n�oJhl��U���������������&�X�u�ۣ"�յ���l�a�Y��2H�4�1���s4zS@�x���s���ǐ�$pܥuyj���%�W����f�UU$Dܽ�>4�߱#�>#lY�i �d�8`��X��aمR�|�!eBQ>Ϧ��ύ�JblTi��R=�Jh���ץ4
�W�y^p�M9WE)DԢ����`$�(~{�E����Ӯ�e�j̻�ņpMudU��n2�by�r�=>�)�s�'�"v�F�Y�<�Hc�C@�ҚW��:���oJh[c��fB�t+�4�]��r�"G��$yޔ�;�����$dq��zS@��4�ڴ
�W�\�vı�Ҭ��˥y���r�\R=���d�	����ɱ��(* �F0@ [
��lh 	O���9��~��@����+��T�/1,xh���^�@����oJh=,J�J��I�D"��c�gj����O5�*��6�8��K�c
���3���W��=�)�[Қ��4)��Pi���mH�oJo�$}��{女U��+�a�udcłk�4������r�(���8���՘��#X��$��u�4
�W�u�Mޔ�*�������@��z^��-�M ��i&�"�`"��{'Ke�횒KS�IY1�|_�)��DOK�=T�9��z`��rk�%�
�dڐJm^8�tn��$S�^��ONb���Z��ɸ����d�[mݤ��h��.�ۉi��v3���=�<�FNb1m{>-����]���'�ir��J.���Aʅ��ǰ>��{6���甠q���$�؅��Kە�ݠ�.uf�@���[[��=�i.z[�ў�rfk��`�T~Z��L�]a��4�m��a5��Ӊ4h���˥��]��Þ��%�颐�0#X��9�{��4zS@5빅	d����?���V�s*���I�G��h}gƀu�4
�W�u��"G�WW��X^bX
��/�@��z^��-}V�}(�c�x��y�@��z^��-}V���$㙠|�
Wb�V�Z��]���:���k��Y�Uz� ��;������z�.��_Z8�v~�^�����u�^ڗ�3��CF�^��u�l1˞;	٣�{��`�w�9�u�Hkw���d�7IR�J*���z�-D4�B�N���1=��}C@}�3@i��,���b�rh{k�:����%���@/��w�+� �ĔRH��)�{���Y�x�����X���'�'!�z����+��x����zS@��V�&�<�1�'l��A�����烡�����9�u�B0��i1<q�L"���@:����^�ץ>���]~z�|(�1��)&���נu�M��W�z���LO��M5�q�zS@�{���<��w�No�<@���BK��"T]�%���krN�߽��s��~1:�l&�r�ޯ@:����w��a�}$�UK.��T�Z�n= ��h/mz^��=^�z��݋�����e=�7�v�\c���q��O[-�նxN�۷6�����a����@�{k�:��������f�{���0�1%�=�Jo�����~���^�}1�qcCK$��t�0�>_uހu���_.�z�!�^�l�����)���?�/o��vwެ���
P�,��H�%$��� J��Q-�,!B�Iծffy�y}���F�H�X�Cq�h��Xwm�g�� �f����g��;Ed&�10p\���݊&�ܽ���9v��&,�M��h�Z y��ww�]nO�4�#q���nh�z����<^��9�0��ƀM!9��ޯ@�e4������׫1G�KT�Z�w��>�f��|��)(���9u�����F�0Y ��n���@}ok@�}�z�s�9��#x����E$�@�n�����/[h�9=n������ZJ�"b�Hm���yۓw2K+\�F����}��u&ӫӛk��/����8v�<�[���(l�u�6@���Z��^v4�]nZ�sˎ\*^r��*��Z��n�)3�7&&厳�`,���;����9���/��5�T��ئ������fE�jČ#[7J#۰�Wo"[��:j�U��u���r���l�!5���ݻ<DZ�MkSY�j拖f�f�x��Ȩ<�w�����߯ݗ��*���K`��<p��rJ9�k]��x�9��v�]��W��n;<�$���p����^��x������/u6cc�b`���z�.��^�z����W�J�Ʃ�Cq�����נ^�s@�{����h��5pCI�8���3�Q�����z��F����K�>w_�O�ƚ0M�9��ޯ@�e�@������ �脽����%G����ݹv�U��@���;?���v�;�D�7;/�C �̱�Ov���o���v����wt���y�˺�ۍ5��1�ۚ&䜿w��8 0B
#WO��R���!EAg��,��Ӏ=vџ�L��S�@U�	R1ff^��Z�_U�^��x�W�w�5��n����}V�zˆ��^����ަ�x�"�܋@�e�@�^�@�n�޾�@��ŎaW��`�q������މH챜��k�%��Ë��nVu��u��1]��~�������`��8�m{KE4�Z$bl��H���jď9�Z�.�����2��F	�'3@�k\�]�`�'f��##!EEUH/��!�4����`0!|?���\d������T >�	�FS����#��(s�g������I1��I	BRP�HZ~hM��������o��c@�V�F,`B2�Q�����@��Țf�����@��Ǉˉ����5�p �Μa�c�y� �BU�!X����F��� $��(u]�X@#雺4L��C m�^�5�>b%#U��"E"1RP�R����C�b}�,F �Bw�k��"��p�0���$%��Y%8��"w�����f~��-HE�E᫰!a$>:0$H������B�hʐ��,"�h�>O��_��? uY�s�
i����R���!��P4 �"��@���L^�D!b�*o}_rC_�ŀw�Ւ��$]J�4�]�М�seɹz�{Z����r��ܒ6��c��	�4uz����}V��e�@��2��Ӟ��n�od���![�G��9�tQ5�͞�mԳ�.�@��-�O�:�ŀsk\���=��~��*�� �GNf��>�@��rw]`m��DDD)��~2�*����@����u�����}V�{J6�E���I0�;��:�����~��	A#�PJ� B2H4��B � F�%� ��A�Z�l�"��#�u�\�����9WW���Q�I|e�k�UeݘZř�[x�mk�u�F su���<��ۏ��&�ݲֹ�g�0��^#O����V�τ�g���xg��v�t�7a@n����@?>���vI��|�{3y�k&�n-�ˆ����ă��h�mh�}kg9U�q#����eق�1��h��4m������ˆ���X��j!��7$��S�����~�u�F su� �*���b��I��<��h�\4�����`I��N��U�oͻ>��\���p��h4��Mt�J����:l��n��fA��Q�Z�oK<�Ʀ�/�
�snW8��"Ocy����cMm��6Lmڃe�Ngv���Mi�9�^�Cv3F���ng�2b鵆�������.b(����i��Yv�E�$Y:^.��Gi��7�i�q��&��e{e�=T>qۗ�͹��bUq\����75Mh֬-˯���_ |��������[\x�^Ó��ȭers�:f%�t�K��]�ݐ�\�����?[o���� ���w49�Z�Q7�АHr5	&����w4��Z�\7�����|65�1�AƤz�mh��֒�T��%�9z�q��ʘ�$�'3@�_U�[e�@�^�@���ε��Q�
,15qh�p�<W��-�s@�_U�{��	W�6,�bd`9�%Y&["J��M�P��&ٛ��t��-k���'��.�s1����@�^�@����}V�m��Er'"nK"�G�[n��q���TG�ڊ�����}t��F��>��=:VK���c��� ���@�ˆ��^�m��{ĸ�,A&5"�-��x�W�[n��>�@�\����$hC�qI0�U�=�w4��Z��;d�K�F^$ee/Ҿ#7L�Q-n{I�ۮx���� ��Y�R���\��1�AƤ~��}��w���-��x�W�y�q��ˉ�l��w���-��x�W�[n��ďl�fb�0Qa��ۋ@�ˆ��^����,��P��	MO��ŀwi�p^�l�,s�M�4��m��;��h�p�/tW"���IV,���ok@�q�_��d�@��u��ʈF�,J~p�8�o�l�Ȕ�˭��qF��!���M�i�on3���ЇK"����_U�[e�@�{��۹�{���Ȁ� ��h�ʴO[��x���ϔr@kǨ�S�Q���8�ȴW}��-빠{��_eZ���lj�cdqǠW��ֹ��Np%B�*N���?��x�rk��7$�y��L�x�-$�W��~��ց�I���ˮ^��n���hb�⑶�dMŀ����s�n3�)�y,t����J����X��#�����XbiF���w>Z�ޯ@���篪�;/U�(,@��bi)�h���x�v�� �js�J"dm��$� ��$�mǠ}��s@���i��E�|���:�ىe�#b�Nf�篪�-��x���m��=�	q�yD1H�l�h.���`�k���1�(MBn��p��v�eh��S3\�q%�c��vjݻt�/c���;�%ڸ˹M�ɜ���{w��( �m��f&�y}�d��������'<��\����!hF9�v�c/��۷�t��jƈ�m�b�m��ǍL��a�FvKngiٛ�	ڱ�;gŇn�\����:p�m"<��e��Sp���/#[k�6��K�3L�&MҲ:;)�Y���Ý�ϻ�����=���� ?}��\˭f�d��u�&�dɞٖYL�I=,�۶�v1���qi�Ď1��NAp��$��>V�=�w4=}V�m��wO�lk�,m6BGz�}��篪�-��x���(c�?yq0X�'3@���h�ti*�/�\�I6��7{�K.�X��ҍŠ[e�@�{��۹�{����l�,�bi70�<^�Xm��;��8n�0D(J'����Ӥ:I}:��淤�/k�$���v:�]����+���r�4[4�۪����$�k@��������~@}�3@�c���D��q,R!9����p��g�kRC�+��*%E�H���T]��+RT/�E1}��� ߟ�@����px�!#	�Zn�0��xm��9��8�R��N�`8D�a�{�h۹�{��l�h��Q��	4�!�� m�X{Z� m�F s�� r*J��C�~D�A#"���j�Bcӓ�(e���T㴏{cz�I�Mx�m��vs�g��OӀ6� 9�� m�X:�٘��#X�5qh�p�=�h۹�{����l�,s�UV� �[���a)B��P�"1
S��+w+y���]�;���7$���"F)�X�rh۹�{��l�h��4.:�&�ıH��h����.���w4-YVj���� @����J+׎X[u%�m���M���;es�۴�k�29v^�=;kH�LjE�[e�@<�٠[n�ﯪ��+�����N)&��v&F���;��8n�0��QSA&�y�rh۹�{���+l�4�m�����i�Nf��J"��~����ηx�DB�S	8����,�c������S%UW8n�0�n��ŀw��p��ؼ���e��Q����pU�j�m��\{p�����s�v��6����J�lss�р�w�6�,��s�6� ޻q�2,B�1%�7&�m���f${�ŠI2Q���͉��ɆbY�j����>�>4l�h���-�k@��n�����b�xhNqI�b�>]~z��hޔ�C���̢��x�2����w�)�W9ʒO����zjI��~�]�?�A_��A_�� ����AZ����DU��EW�* �����/����
�H**B
�@��*��*  �@R
�UH*P��`�@H*b*��
� �H
���"*
 Ƞ H��H�� �@������D �D��
�
� *b�F
�`�B
 �*� �H
���H*��E��*R
�@ *
���"�E��D �A�"�"�""� ��"�
�"� �A��F"� �� ��D*H
�X�
�D��@`�B���H* * *`�E��DX
�QH*T`*T"**
��"���*
����A_���*����DU� ��EW��A_�QU�DU��EW�TA_�U~QU�1AY&SY�)s��ـpP��3'� an�       �   �    ��  Q� � Ȓ	R IT
(�P   ��� @H�" � P�    @*R  !   0�PR� 
 U� +���ͽj\��&���-�o �^�qoZ�6�맣�[nO]Ox@<������ v�uW����} ޕ2z�\ھ�����ɧ�� ,t;���"}t�}���� �   <  (  R�X S�'��r�[Ө��ʽ� 4wϩsoZz�M\Z]n,�. �Wsuv�-����rU�)�7��_/��ک�X��כK�.T�x ����^������}��3��� �P �PQ)� 4s����ק��P3��J:DiJQ� ��;���� ��QL���7��:{4��l��JY`� ��R�Y`� �4�� �A�FvP� 0�G X�Mu��P;�Ҁ14 \r�J @��� ٠ҌJ�K���ru/����� ��ũӖ���x�u��R�@ҽ�'��� M�i��n�y�N�^ۓ������x�]�o�W{� >�Jͩ���6��n��<��M����J � ,
-���[�����yڽ��ͩ{{Ş��� {�����R�o;��O{o6�{p ���}*���W�/  /]���������(�J�o�ܷ�w6�w+������.����m{^,�W6�V㺕x   ���m��T�F�"������JQ�  ���R�=Hd�	����R�<�T�  ��*m�JR   DPLR�" <S���_����|��c���r��q��` EW��_� *� ES��*�� ���UV*�������P���0i�&��gP�����M���i`Q�H�bA�c�?���f���>�s��e�� �ć� *ap����%!��ٔ��	C@#\� U�	1�%L�$���O�� �9�6f2:`A���pi�WM"Q���CI
r�H0�M�.�%�`@�(Š`2F��s���
9�HS!��a�p����s�SPa�}�N��M��S���؅�U�D�#@�`@��`Q~�M80d$���|��"2 ��BI!$`��:�6�+*AZ1�H��M�o>>oF�!�l�jE*�2��2i�, aˈ��I	zM���X�sZn}	1��K�n&f�0�t�󈔮 !q���X\+��\P�V0i�|e�BG��3��
����́��M6*����`��4�L�k;>:.���Tk�%CD.�P 0�W�=:JbZe5$�2�1&�7];�	1�m4��8D*8��#�a�	��i�}�h`X4�$� �H���ҕ0�2h�����
E
� ��؟v!��Z1jD(���+!�i$��5�fmbgV餒h �B��\N�ٚ�B�����
I�Q��#e"F�Q̄�+*�$'�܎��A�+aLIA��` � 2 	P�L?:9��������sgP��0"Up�����^��4��	0�B]Hj�N�U��!q3a
:�gU�h a��:����D�+��"	9�1��&�"Upd��S0"�4H!3��o��nRA\E��432D �p,&����0)��Bs"G,��-�����5��@6��))�#�D"�b"B a2h�2�L;��y!хpf1J�a)�S m��J�P�@jrp `$�3.���u\����ٙ�&�-�5i�ݘ����	�.B�����I���_V}�$�@�x�	�Z$���`�G�㖕_�.��Bf�Ʉ"� HD�!W���B	�bȐ���@$]�,&����X#~�I��0v(aˣi�d_�d0u!��H�%d��[P�WfMJcSQ���fq&~��	��Na��?D(���S	&1�i�#$eHWI
H�$#@�A#,Ę
����S]��� `���rD�B(�G�d���jB� ���V3�w20*`ɗ�-��@�
Ƹk����H��4�a�j�2m�0)�&��\�B��K�f@�>b��50d�ٟ��>��9��ϓN뿟�b(`�0�L8S`4`�XBY�P�$$�JrW
L�A�@! �Q���	��P1S,�D�(���Sn S���HK2oX�c>.�h@0@�@!���f9�r�gy٨�Ncq1�� "��p��L[�lY*.��>��%b�d�3�D�VL	�h�1����hHP�� 1�Dr��3,ab8��aF!a #!rh!��l�N�>��Dh�h� B���đ. Y1)�@0���|N�Hs���⑐"@,�dX@��L��}u��$ RP�ɜd�+�	˭�f��Gj6bS�vR��7]�b$Jc!�m��ư�����l���1��d����]䔎BH�bS�Z`�"�W�A�"G(����EQKiȆ��?����B�aL\v���B!q��
`2d���H�j��$��p��"�:�g[Ѩ�)���A��J��D+��C�0B�F�}�D2,B��ɤ�3���L��T#H+a�@JB#��U0)h! ����*!�.w��逍�Ͱ��l���7W��Ԙ�.���ę�	P����"�H� ��U�Ɲ޳�6G��������.���ނ�.+j^ %��H%H��~��a����5x���ĚHĕ��&����!�C
�r���'��4B��.���p��3	'y�&#�%�.y>Ӓ1���~6��.2O��u�ID��	�>& ɢ7`s|�+X<�)�$��!9�A�:��Go<a-vSe���\:��Z��$I�(htv����Cd�5������SK���g���Ci�F����c8�B��N�����P��N�K�#Vp#�a�f��ư�M&����3��4ټ~x}�D36])��3��gp6���q�j`@ɢ2S	�_l�w�S}D��5�f̤��X�,�����	"��2k�I9KČ�Ø�F�!U%$��r9	��J�8 Y�q$ޠe�}'^9�vMg0��l΍�r93�w`C*B���ٙ�����uApuU��/V/���b��U�ʯ�/�V�߸�$}_��ʯ��4��@��F��}��f6�~)DtC,FI�J�V��B`����Tb2XVA
�;4G$X1,.��*F6�@�)��]5��$�Sk8�8���΄	��9#�~,�e���X��sN�BBFI�͘-0�p���O�!38�,ÕH�`I�M��\��B����@�K�V&(J��9�|��9��gF'�~W>���hO�DEx��&_�pn�tٮ%���hA�"��qy1�+}�y��2LgL�7�![*�i��ɜ�
A�B����R�u�o;ɗ��e��vl��:'�)�&��.5�F�,�W�H�*���
!0bB9%��|�& �&��!�LJc��:t@�SH��%@�H���\��)���e0�Ԏ�&����ep��h0�M	��C�B�28�B4�4�i�nv|d2!� D�JH��## �$	(�`H$[�X���a駦Σ�l�9po' � �cN��B�2���:�Ǝ$��) �H0 �`�E��%�W��IC@B,@I�X�5�]� F@���d:��X��)7��K��k�g{�g1���Y~ε�`��!jF�b�2k�WA�%�)�섌�̥�oB|kd>����H1!�����3�4h!BS,���K�\$[w��]]H|G�r��P�М�a$r�8 +�2k&Cd>���	�F�D$j�����L�8Ԓ���.1�0��Ұ��0G&f��9���w��B)!a�W
�!	7!e�3���Ak��,,���kI�/�^uR��&:c�����@,X�����C	�HBf���!u�\�0��BB�B�H���ǃ��x&��b�sF�7)��X�!H�)�{\:���[7�D5##&̥0CIL+���A�n@íGlI@�O�pl�)�`��&��B�&��e��
B��N~	p�4M�(K��:e0g�d���)��Y�*3�B�B"�H�8�&��D��!�A�>!���6��a�F�	�`�4��� ���      �h    h      Hm�       �` m�    @ 6�            �n�         �   �`   lp        I�6ۂ���-� �5���\�[@8[N	r,ʊv�\�6Z �h Z~���  km�   f
UZ�z�U�=���(��<���O+���ma���I[m&�n�ж�X`s�/��ڰvE�I6��n�*�m�4�T��5ЂY�y8�0����-��jUu���;D铗Y�dq#�Z��n���}~��:W4���bv�SQ�������	l��va�""Z�VZU����\��Y�m���)VWl1ʭUT���u�g�(nk-���b�l�Yb�(�͙���Z�6U�Dk��Iq��X����m������Ij��d�������GMm�%Uڹ6��W���ˎ�fg-/=W@�	VJ��
ڲ�Ͷ�m[\��I���j�+�p+j$pl�.�[<�ʉPm�m�P:W���[�$:@-T ګ�
�V`��vড়�N�nb��.Qy�ڪ� ��m��ij0p �D�]a��������  �n 6�����  -�^� C�[G  �j@m�m��]��Ƶ�9�ך��'n��d���ʒ�nE�`E�m�ͅV���lp��v� ���� 7c�	�@N����*XN�
���V���Չ'Q�IK[i0   $W( � �
l]mT�*�r�VLl-d��n�u� $-� ��Q�Vԋƪ��8�nm�p@���:b��ڐp$!��\#�-�۰8KZݖ��$�m���R�0m'V� ԆN��U[Ue��P8�eِ��%#�U���@�zλ�T��m�  ��i�.��YAm��I���z�~��m~���]{$� I�G� 4Y�I�ސK=vۀ�U�+����j����n	0qz�n�.���2�m&�h$ s�f���a�n����7Z��hhQ���\�hY[����]��  r�/YB�ۭ�j�,�_N�Fc���%3���duR�	�̜���p�	���n'd�v馉�ղ@F��΀��Wh���5��\ k�`lH    ݶ[m��]�[M�+pV�`r�]k�A�E[l6Z�5��H�$%� �l� �\���Z�'P#mrK�4�-��  ��,l�wm�@ � ,;I��p H�U�$��߀'�'I�p�6��l�irP-�� � �`��   5�k�I���o� l��.� ۶i2��mHr�  8�n��m����� 8r@��H��m     m���I�E � 	� �m�      �   �nm   6�6�  k���հ ��   m�   -�kd� �����@� 	Ԁ	 �%   lm&�I�� 	$u�^����pl���  �� j�[Cm�l��    m����mf����[l-�q��	   Ӏ  l�*�J�6U��MMu   �   ]��^ăm��A���t�l�m���M�UTf��;U*�  l:��ky&i�,s�
�T��N��ڪ��@��[$t[U�;/�-�j�v�]����e[���j�nuLZ�Mٝ��2��R�A�U\��9ش�Y1+�e�h
�8%`��<��J�P   ��m�֤6���V��$$ ݦ�kM� 8  ��&�v�ِ)I8ݦ�t�l  ���Y� $�R�m ��/^����l�%��m�   -�kH6[@�9�m�p�k[@7&��˻� 8��   �m�K:[�l �$�:˶  )�^Vm�Zq$�6��d��m��nݶU��� �vm�d� l�A%�mo\��-F�I�` H���ƮͶm[@msl�n��m�mRl�ձ�- �	  ĉ4�FhM\��JA[kK6W �v�[@ [E��Kk��kh ,�d�����m�d�m�$ ���mM%�aÁ�$�YAmmul�6� �� 9�W�I�WM����q�<�KP�ixܛ,C��7"�d��	��p �&�}�M��Z)� ��I�����!סR�h�t�Zm&8��N���*�K̼��[m8�$Y,���i6���K�)i���
�'�|�#����7l8[]�յWT��ݡ]�T�A��N��*�W�j���cC�H\��%^�V�Nkj5M�Uuu�����$�� �n5�;�ʹe��0ɐ8^GWX0jY�Fz� 5TP�����"m�e<�9�hy�wf몪�[���pi��K�]�6�m�m��JI���9tٶ�m�mmUm�f���̜'�յUe%@QT����l��	���`���ݶp-���A&���u�n�l H��a����j��Ԗݶ˦�L��d��`�8  H UT�*���Z^���lq��� lkV�Y)��� p� ���@-� �e��V�   $�m�   �l[Am����H7Y� ���� �Tu���'V�� �kg�ە��A�]"��@p��>$�� ��P8M�6�I�h8��כH����  ��Rl-��     ����K��[V�۰8v� 8 I��v�m�HkM�[�e���-�/  h[d �� m�� �����v6ٻl�d�k ��ҭ���PP��\-�vݫf[|p-�I0 6��i0~7��*@6�m	 -��ו��c��h���lp 5<�`3�UVvųʲE��WJ�nI��r��+c�<�6�R�����SH�
����e檼�y�5�i��Er�cq��[p�g�_��u� H�H>��M;O�R�Rػ`  6ۀ�]n6�-�����ѽl�  � �im    �� ���ٶ  �` -�k;Q&�I$�ۨ pH88-�n��I sZ����8-��d�� l�R�p   �p          m�`��la�� @ 	�  �dۖ� ��m��@W-����Y��l  �� �   ��.��� ��6��m��vm�۰j��q���    $�r�m[�6��Em��[��	6ZZl !�$ͳluq;/]���m�v��l��4�[I�6Y:�� �� ������    -�d�$  �V��p[��|�mzf	�����Hm�	  -�6텴����5�R��l H��k3�mH��U�5��Ͱ�17f�rm"@ kֶ��$���6Ā$ �p    �  6رͶ� rE���i� 	-�l*�ڶ��:�R.U�t ��ݪ�[�ڪ�r+J�e��������m �Y� ��t�m �qm�0	��   sm��$p���� �-�I�^��$!"ہ���,�h:��&���N 	���KW:تt*��j^�`6�4�[P��Z_U�Ȯ�T�v�-�Tڱ��e�Yʰ[[�q5uѫv�-�������"�.��U�a���5�TmT�rUV���J�)Z�W8l�����f� �^� m-�Hm�9�� �p]Wv� ����(���  �m� 6�n@  JV���p�I    m�� l   Khm[  I&ձ [���Հm� �'1�Ͷ�N����`q�m�6�[@�6�l��� ��`[�	@ m:fm�[ ��`   �   ��v�   �3�d �u�� �  ��6�     �H2)$Ҷ�l��:M�l 6� �am�� � V���K��X
��P2���j����U��8�m\`����T��` h/Z   ���/Z  �kCv�i��Ls�E �5� 6�l�,�K�Z��������B���_[\�ۓ��UX�s�I;5mI�U ��Q�l ����غ�m�[@ հ  8��-�[@ 8��� � �� p�        �ŵ�Ŵ [@ 6�BF?���{��w���� !B �"�A�BA?��()�j��E�?�9G�s�i@`	�B��<:#�~ 4� @�e
�Eb�� �o;US��40�����.Q@����TS�@> ��;�L*@�A:�tm�X��@���ʂ�QM�pU�QJ@�U2(	����P6�*2��CfAN'`	�6q(<�XX�(]��D~ �S`���PS�b�x)�!�HXA`� ��$# A"��h6���@d�N���"�N��� N��ࠆB@������|��L#�&��؈]
o���iD�	��mUPخ@*�:( І��Qb;8S����U��=6"&C΢�� (E>q�> �~0:N�ꠅ�`!�6��h �
�#�"#ү�2
��B"0F��?<8�!�3HU1S���Q_��\��vK��ET� ��t��H�$H��m��9��p EWB?�S�@b�� �Dd"��E��j���1�c�s��<���l�$��  Ik��m�YE���HHL�g�k��� ��UESەݶ-�hL3�JY-�a�8'��S�����Qp�J����(i1a�N���(q�ն���M�Ʒq׶�^iK=�d���s�Ѷ�t�vv���&�h�]V3vwnc����i��ͫ�����pf�Bz�V�N:���'�çHb��^RƓg Jw8�E��$����9[�;.��n,�G��;��m@�䨀�ت̀=��
]���k�;�/-���[)��n�[��3�U��d��׶���n��U2�#�+˹:�Z�۰['i&7[֥���U�8��v3�
�V(h=�m�e�IPъ]��C�V�L�/`���\4SŁqѻFLup�\�
,�÷k*kJ���\�|+t�ol7Iӌp�u�]�z��0����\�i.3�N�һ5T�/���m�c��zA�֗�H�������vJ����d^;>�iը�L�$7A���^+�9�Q�3��pg��ۙV܋��/<�u���:���v��z#�ى�M��Y�ڒ�bR#CV֧��X8m�Ed��	�5#�nА�b1�-d�.ͰM@U\���J�)E.���iۮݺ����i���LsPe�;&�i����Q��Ƽ۶ܲ!B�6Ύ�jE����׸�ssN�ܶ�"� +ѧ:'��q��]����B0cV�*�J��Y�*�HU�Sj�S*ʵ�xydɸǀ�mv�aT����L����3�Um�7��]������F��,���&�J1��L[��1[��,Ԩ
�R�X�
��"5܇N�ʩ\��U8���$΅�g2fۃ�tUn�[R�.�u� �kn	&�M�е1��s ՌUl��4-�m:��eZ���ե���.�T�T��gcs���-�f�gA�75 +v�K�IN^Xԃd2M�R��� �d�q*"�P�"��<dE*�c D��SBm�;T �)6����~:(Tf��e�4��/¦�Mf��560ӹ��4���n�q�s��6��{qΒKA��1��2���ԥU'i!��;Y$�X��TReK۶z�aT�4,�"j\����q����8�v�a�������z7*���l�taSf[U�olW;(��8֝����͠��u�b����^{v��Gc$H�v��aˢ�n�����򠦜���Բ�K�I�b�Zb⸐}��ܜ�&��'q���p(���9	 ����ov���U��/���;��,|m#�U��������ڽ�����B���v��� ~�ۀ}�dZ�NJ' �NSv��� ��H�M@{� <���j���[-X~���ۻP�EH'��$�H�b2���77C��@�j�%�@6�nb�?=��[�KcE��UB�YH�G�n�p��'��ː�hɶ��6r�ϓ����W�e����R7 qR ߻� �t�ͮJJ����¬~�����1� pom�������?}��`�V��l� qR �����֩�*@}���{+Wj�Uڰ~���ۭRs���� ��ɛ��Yw�����n�=�Z��Q�T�m�Hsۀyq=�����]T�!7lt���{5���R�q;���ΓA\�1�ճѓ�p8��㉧-u~�o�`�w w���?}��`ou�
�W,��Yj�qR |�=�Z�����b2��G[A�ʰ�wn��׋� �9�(��j��lD��4#� =Gﻏ��P;�w�7���Sl�T�#����j��*@6� ��@u3'鷙�m��n鹗���qR� �n��׋ �\]�^^q~t��"@X�L%���۷L�kth���ݺm�5���917!a�JIUV��_���b��ݸ�^,��q`vv96Y��Q��i >sP�-R��H�T��t�)d:룍�p�n�X�������q`~���b�$NWc�0�UM+�Ձ��ՀgqՃ�Ӑ���֌3�	�DЅ�s륀~�|�ʅa+�V�,�`�w gqՁ�[�V��b!B��H�����u��ve�gm{ �ӭY�u�O�7Gf�œ��f��}�\��9�j�27t^����ڰ>x�zG���`u��~�6�eN�9n��׋ ���H�T�9��M+%��f�[�ne� =T�m�H��Ij�~��>RJ��Gj�o���X ��@{��HG 9�<˙������2�j��gqՁ�Gsv~_�{j�s��I6���)DH,T%`��IHU*@�jD��k�
)�B���L  ���8P�n�w��I+x��-�ぽ�oHtdz���+[e�/.�2q��n��<kt۴�;C��e3�.XN�Mal���J� ��;�r�j���:�Q堍�
Y%��\�nX��qK�v������ў�����W�nqͰk��	�7d�s'&�� �Ϫ�Զ�ܧm�T=��*ܺ#XwuDr����#���q�H�;J졊������b�)8-!Ul/���%�l��tƱ�׎�����^��8xy���yBś)d:룍�z����?ow��q`~���b���`�+���(�{j�=�猵`o��ʅa,�W`K-X{�ŀ�5�������������"NO)Xl(��Ǐj���-X<v��{���7���Sl�T�#���������� >sPT���@�n9�Sѻ��헭7f��#v��^��ub�Md��=s�s	f5n�����R� �oް�¤�o�"���Z��X{�ł\�:�(��T:�ML�%�p�����ō����5��a\�����@���������� �;I��(��W#��y7����;��n*@��L��+3,��q�v����� ���|� ߷� ?ot���ѸI�WS��>�m�V�A��]M���9��:;c��K�Q犆n�a�������Hm�@����p��ŀ~���&�RF�M�,��:�ID�w^�`w^ڰ2s,ɼ֞چ첫Y� ?oV���qd�� )��zy˝���Ƥ����˦�9���5l�Un�{ �9�������.�v�ʪ�Gj�:��� ��ۀ��n�{����vR�Yd���n-Ps�Q���j���l ��T�$N(^Z�-m;�q�$yl�Er����~�� ��[p��ŀu�ݘ��m�"��]j����'W��)���Հ���3����;����9]�8����o�`��@����jt��������V�ȗ&�� o����Յv!$BP%
%.uӵ`co����U�~���w7�5 {�5��_�ـ��6AE�[!KAȭ��s}��y���|�7�=�sk���p^��WGdμ�T��[a�����~��,�����ݸ�5Q͕���e����y��(�E"#�9��ﱠ�}p�ۮ���F��ʪ�e���s�5 {��@z8��b�m��d�m;,��ݸ�Z����]W��V�	��ܻܳ,�+o2�u�� =T�v����V�B�\����rSNyEU �Mf3n��U捎������EӺJn��[��d���Iz-�����]\����.6ꑟsBLM�x��o	�e6�2����>~=�h���b�:-�BFՃ���<�y����b�Uts�V
� �a�`a'���ۍ�F����[�W�����C�D���c6z�pJ;�i	6���Pq7e�:gd�P��x�k�������{��xC�_�����Ѯ�\��ܛN5]������۫�y��ݍ]6Q�r�6D9k��w��,��ـ��p�n�X���,r��	e� ���Ij��*@z9�"9*qB��Y���p�n�Xs����ŀk���>f���vKT�y���9j��*@u�1 6�>�Nl�8�u�ku`�w���S�>� I>���T��(1m���..�Wl[1LW63/Pu8��t<;�)nd�w�gX��^f��m�@������W�Xt��H	2�a�db��FӲ� ��ۋ�I!( BJTD��e��nՁ�x�`j�i�UG+�W	-�;�tŀyȩ�� ۚ��2�fe]��fP^i����R�9��5 �� ��]�E��Y\�-�`=��RIo7w� ��j�m�V�+�oo�����Uv&�f�������G�rzX�kok��:H0;:�jLXU���λ<�v5���>���� $�R�9�3xi����-��f߷V,�9�&�{�ŀu�}0{�0�M�sei���R&�+��X���vv~�P�&v�0)F9!:�EҨn*@"��@��!�g[�@1S@��$$�AS �� 6�b,4T>5��1��cJ M�`D�9���I��)���ƻrWJ@�F��sb�!�\��D*����(�ߔ�ʲAC�S �QnDp�A@0�8q�h�Q�OQ�@J��:�Tp
q(��9�{?�Dݓ�{�F��l�����[�^H��`~����`������KVS���V�)����r�����@���vG> ;��\s=���I..vy��`���Ii,a���F�;v�W�[��[�dлc�3\�ݳjj���u��r��{}�b�?�����_��6ow����^RDܱ6��`w^ڿ(I/G8{y��>P�M{�=�yb�\���z����,�W K-X$�N�{6�D%/��nn�V���wf5
�]C����wn �ڵ`|�ڰ�԰��D$�1B�X����t��u����}g��D��%��� ߻�,���0����t���fW,�	�dN	�S�u�;f�J���qY�֭q�g�x�{V�ùvE ����']�`{ݸ�w^�{� ߻�,Wyիm�ʯ$�3u9h	q�@NpT�$sP؛��ꊌ���J�{ݘ��1`�v���x���v��`����f�wLX�ݸy�l�<������v?E�$c��� v��?$���j��ǳ�G�;��}'b|���
;��v�w�ߝ��۷�]x6Y6�5�C�eqy��M=)�d�,�3m��kn��`(0vh��^�$������b
	�1���Bp�S����s�z@w� �t��n�π�3�MG`��n5{[�g)�eڭ-٧X��P6���X�s/e:�\N^����1���J�vP� b���#}��.'n܇se�����m�!۱ۑ�Ō��s�֋� ��B�\]����߹��B�5Zx��X[&�f�ܶ��w=�9kp��ۜ�j{:����n'"+C2Lff����K@K�bt�� I%�?wvaP���q�^�wf:JT�$�P㖀��B��sj�s7k7t��@N�� 	$�x�#�ـ}��'6q�붢¬ �٨��@K�bs����ԤV����ۀogu��v`��ŀ�� �ψ1��[D��["��#{��ɎE'�
��qm�C퓆��h�D���2��\���v`��ŀ���~a��j��Φ�q�Em��~mZ���P�(IZ�QTwj���\�{�3�l��輤�v�0���� {�V�c�6""!L���}
>���V�{��V9c��[m�7���rL@N�� $�������Fa[�n��ܓ� $�\��罜��KcE�ƪ��r��tyv�k�U�M��|�����9x��.$K<M�fn�n雸�|� 9&�:㘀owf�E��l(䃮ڋ
���Pq�@;�b���ԤV��^X��=���wf,�|c�L�ȎQ1�s}�5$�w�Τ�؛��c������0�ݘ~�j�9���ȴ��ܲ�
��f߻�,�$��޿����`{�0=�����Y\�q��
����F�F�ެ.�<����d�vz2b�y{UC	�U�}�\�ـu���;�tŀn��+��Y[�V�p��偒�偝mZ�m��P�d���8*�!l� ��z`�ub��q$�7���:����ׯH��9d�r��Ur�aBR�u|���X���R�H	 A s�g������<z/Q9�Q�]�J��w�c9�y�:��u�k �\�R����JY�XEJ�ܯm��v�gh��K�t^�8��d�p����w۩�J�-q�~_�������;����/��plM����Elc�`=����K�5��Հk����|�21�l�TV1X(�`�ub���p��f����>��-Q�R��)�j�@��\sq�@>�� <��+��Y[�V�p��f��g�y�7U� ηV ���!"|���y�.��7��������fgsn&;i��FsN��a�lQB4��c@X��ʵ�&q�N�p�T�rv.�z�aƹ���MSrck[EK��V7��1;!'g.M��lttMt<�[����^�3VS8��nP;:����a��M+�t�,=[i�6���q�.��z��=���n�E�n�H��㯲�S}eÜ1�yn5��=������ﺸh,B\�\�2��=�wU��Z�O�]h�ſ���ݻ�r�l��[.Φ��l��,�jՀg[��Hd��X���D��%�[	,�;���g��ĒR>.rH��������ئ6��ov~��s`��rH:�uXcm�߷o�Ͷ�EX���9�����)`���ߧ�R�Tq��R8�6�^�)����ݟ�6�f��cm�߷o�ͷ�z�:�+R�1�T��M��ߛo�ud1����i��m����o�n�Ͷ�N:����gm�uܱ����C�<��#���ӣ�Wj��,��Ec��Ig�ͷٺ��o�ni��m����o����m���X���0ą�L�j�o>�{w���6�`��r^*�o���ƭ��s����O���������`{QG�����)����ݟ�?$�$��,�6���y���MلMB�䤁-v�m����6����cm������ߗ�~��q���y���%NY-R�ܯ�����Ym���߼~��߶��m���u���z����>���sLv6��7l�3�ݺٶ�vd�^���XT�t%�����q|�qv�s��o��i��m������]���}~~�cm���yy~q��RB�~��o{v��DB�^UU2�{���3>�x�˙����>��#��o�#�*9e�u�^6���7�m��f�j�"�F�P���{�|~��o�}^6��;�6~UEc��9g�Ϳ����>Sm��x������x��$��?~m���(��j@NR�����sOߛo�۞��m��}���m��1Lm����7�$tv;B�&�Q�Eb��M:v�'�H�O/���W����Ȟ��<��}����a�[e>��߶��m��}�~m�{�)��6����6�_�0��X�p%��j����&�ʪ�2��*�wwm�z������ ���?���[�Zi�����X��﹨{�ww͵www�}�}�h��rH:��cm���i��v��=�Զ��y��v�'?:�� @� 2!�1���!!�jHb�`M}�=/�Cm��s��Nڂ�-��Ͷ�EX��謹`��z����]��������A[Mg�ɷJG]#�� ���ewa�{m��[/$�BU�'8�p��YaeSm���~m���������K�o_��cm�s|?9�UU�V
I%��6�gt�g�I/[[��x�����ئ6�{��������,QH��㔰��{�柿6�^�)�����msw����پ1Lm�����j;%���l��ͷٻ���ow�~m���co�I����ߛo�ޘD�,rEdC-����no�wv��V+����{�ww͵vۗ�8�D���� ��,���+a�!��"A��A��p&�)�L�d6$����arbBF!2�"�I	�1$	'�9 ��"Hŀ$D$��Og(`#@���ȑ�0`��H�VTbD%G�$Œ�H$V������S�{����!�TM$"E�S@��0�X�`:�`�b1[(�+�1@�Fn� F"�"0��`A��"��$X�Y��I	�0CG���e+#HD��XF ; FQ�`�	Yg�qA���"�3M1����� �`�E(ŌY��FA�p������B��H1%=ۆ$ ��dfʎ����e��H�`d�LE�aB*��A�"��ۦed�.B��IA9?@� @ D�A�$	!D�$H�HX��oN	r!�F@���Ɣ�@k��b�D�"�2�/z_λm�� ��[d�	�m6��� ����:kmmEh��n��$��q�5��=�N&����u�;��=��=nk�����Cz`���HG8k��˺�s1����@�.֞+,놅%^�t�6N匉����+�[Xq�lZ��l��l��\���=���;[�� El=��Q9���U-��>6���
�K{�"ˣ�9ʐ3��G&�mp;I%�ҁ�sZ��֓O<�[q��kk�1���.9�9���p͢�v!�cg`6r�ul�Q��T�b -UT�3���܋ܠ3�X*��W�pV���<�/"����ۜ�k�æ��RP�8�N{\��D�t�j�����Ę��ͷDUW^t�̀��a�^�M�hm\�A���y�wOj{\�#�����C��S��iF6�U<���s��
�c`�R����Cu�CW���Iu��I�Z�Ƚ�X:m��Ar���J����zB���&x\�+��"J 2�M��;Gm;�2,�-�������n���&�Xs��;<muc����ɒ֫j�����:���Tn�cc�{�"h�m�F�Aj70��b;Y95F���D*ɶ�-0Hia��4� m�BYI��t���Ӳ$�n�H9��mMR�홎jr.	Ѻ%@lǃ�&�cM��U)�;Yvՙ
������ך�`�^E�`����m2�m��U�Yrc�5��*��lm����$�fs�V�%YV���YSpq����9:��xi�45���ڪ���XU����2@�J�t�:jP��~_�j��<��;�4��#;�YV\\<�h�
ds��.:!�o^uS��"Yky�L;K�ٟ6y֡eۓR����*�F�Pu��5����X*�Uv]��}O�!�*�K�,cU�L���US�\��nһt7*`*�Xj�Z�5�yf4�3=t��&HԪ֮g@v۰ 9�vĮ��!�oG_o��	�����6"�G�H�p,d����HN�P]�:3��M3��E�s������\q7�g#���kW���j��`�)ݜ�k-��)�h��Og��;���!Lֻz꬚���.��yM�$�Գ���z�e9��+�xѹwFccc����6�B�PͭC�bب��`8O[Y�(� &�6�w�}������ɉQ��im�يH�K�sk���&J�-؝>��w�]�GLݡc��w�#��g�FI%���Y�ny��-��"��{smPa5��\7$�3�����EX���F��]ݼ�`���ds=뻾�(��rHX툰�cm��柿qqI�{!����}~m���cm���;��Q�-��-v��6�f�Cm��v����qI5�Sm�<y/���z�����Tr���m������6���4����7r�o�n�\����+#��ߛo��b��o������{۵�`����~~ D�"�G�-�i�ɺ5�됯l�Ý�u�n����۫��1���er�sͩ��r�Lm���i��m�������o�ͷ�t�1�����SQ�-�`�9�f�m��{�McJ�@XAB$D"�a0�CGS:��G7޻����ݸ�=�UVf[��0��X䔑�Xcm���_ߛo��V+��q�{�wo$X+���អ���cn[��m��LSm�{�~��}��m�q)&�}~m���O�r;b,*��o���������cm����ߛo��b��o�v~�;J��Wl[1`���eczwU�qd7go�ka��3h�������G��Yk������d1��ǎ��fg'k���^K�S3�����3>�p�� ���q3� �����??yQ���.ff^���fs�����eǼO���UX�`�r[��m����1��w�����B0%u��q﵉�m��ﳽ�oq͋��j((����o����������ͷ�=����o�ݿ�6��g��J�o�{<;�9%��b�~~ �h =����v��m���Wm�{�~��o��;�5]�g$\�gc��&C-�Y�ιK���8G��l9:�an������ǙE��u3�6�{�����ϴ�Wm�{�{������d1���ߓ����cn[��m�i��y)#{���6ߦ�!���w�~������2G���[]�m�<~��{;�o�G��_ߛl�����o�;��~"%�j�m?~m�z�Cm����ݶϻ�۝[Mj��`��������u��������oLk8����8;,1����o�Ͷ}���o���������cm���v4�c%���4#:Ѱ��gW��DOѡw���{\��L#u�I�������������C޲�[��]�ݸ���wr��U���Y�^D�ٍ����?~�?=�)�����׷ ��u�T�,v�D;sD�*@9��\��`���f�5K��"ʰ�ݸ�u�{�*@F�"������������>n]X]���mX<u�%L$�%��I�!읧Ǭ�r�.�V�����ݑr��p���En2�.z+��-�&1���9ל9����N�0�f����/:���=cd��l[u�mcđT�G�n�(+�p"�fGg3�8;d� �p���F��y�c���������]�ڂ�=��`7e�S�|�B�,�&�rӃp=�؞8�i糵[GYNn|�bs����S36bɟʪQ��kR�:�sY�K¸�D��֭ێG8.�`wi�Uέq�g���;oj��;�o�".�F���fV�x�X<u��@���Xh5��"��j�m0��,�a��\ �|�p�n���oT�#��[r�ͤ 㚀<��@8�U�|�M$�դ#�j�%�����=�� ��e*��ڽ��o����@8�T�sP�{p���Q�m,R:������ۖ�u=o'��	���˅^��Y�[-��Ehu��.鵔^�h����5 tw5 ��L��f�5��"Z�0��κȫ Sqe�㗹ԓ�s=��ۦyq..6{t�Kj�9m�7y������@>{��@w>�=�X�VZ�k� ��t�7��0���7����j~f�Gi%UUUw)��9�k��;Vu�0��l{��%�咻iu�;f��6M�-��V
7`�v��8��M��W<�G��wr���D��@�@8���L�i&&�$v*ԎKp�캽��������u��c�V��X�-R�
�J��;��`�n�>.|�Q}���� ?o^����
K��7kh���9��j ��jqs��<`}��ơcrQ�K]� q�@�@8�	�`��������_'�:.�v�ɛ����۶ãZ�:h7C�\��Pqٲ[�#��%qCV�]�n��/�@8�	�`�sp����B����K]�w�Ls� ������V����ͼ������ 8����� ��M�2�⣖���˜��{V׳�`c�e��J!D'��#������oM&Q�c���#�� ��jǰ@N{ 㚀���}�1�����uց��^��Ns�����xvػ@�s=���us]��acw�O�� '=� q�@�@zK�
�����Q%��7��0��� ��{p��L��͌|�G%D�5E�u� �\��R�Q
e�֖���@7$v���cn[�}�j�� =� ��;�B�,7//0���3v�P��9�G5 }�{p$��qw�E�-��Q�V�Q&���k=�ۣ�J䶽˞�^�&z���uSu��d|��%��mY�:�����v9������r%z�QYW\=%�b�Wn�&Mn���$[�6�q��h�[�a�m���n�����;b7*��9�7$)�������q��w4�[A������^#\�(���;X��gD��=����Y�\P�Ֆ�v�2�-Խ��6��T��!T�(�]�����x��<F6�Wl��:��ݦ��l��v��bv��m?���ov��׷ ��t�?wS{�8��8���j ��j�� '=��%�2���b�H� >޽�~ۦ�v�ov��v,MB�-B�����`�������Uv����;޾pU5��UD�S ߻t���V޹u`g]2��Ic4��5K��[�����Ӻ�v<q�BuX��v����ju�zx����$��H��d�+"��������sP�� ��0.�,�� ��ܷ >�^�KV��ĺ����~ˢG�@9��Ы����+sv�r����7j���2��&L{�`�;p�A׫݉�;ʭ�`��L �� �\���Q8�����Rs��,q�i���pq/M�����,~�� �;�3m��|��M�)fpl뛺�X6�`��/0�nۮ�p�u��:������8X�R9-����}��,;_�"!y.��z�{��<R�R+k ��q��H	�`�<����ٞ�g�����+� Ij�=�Ϧ��|�s�M��8��ɗ�1�6�1¤A7���؋"�>�B�tCQ>>j��'�r�"`ÈP�n��q100A��P�9Fgt���ϲ`��SQ�KaǆC�J/��2�s�r��J�N��`�a�@@h ����A�D�'U�e���T>�"P6�AȈA> t!�x��R���r ;D]� �q�q���{����,��I�|�I"�!�ʰ<�w�-�}��*@8��w�Uv�cn[�u���������}j�3�Ձ�����2gT�6J�Urx\n)��8��{Y竎v������뱌��L��W���$���,�}�ŀw\T�I�}Rb΁�Ee��^�{�j�v�T�I�}Rb��`����j�r�e�ʰ�n���0��ذ�}� �|wf�lxnV�f^f��u-��HT��}�v`��bpV�j�E�W�}�*@8���c�h���W[���1q;j����Oq�ty��M�Ǭ���"ܫȝst�xi�u�%QN�Mw���~�R�I�x�Z���|̅��d�+",� ��v`wn� �{����� �����1T1�m�r���B����T�}�Zߣ*�A�䂶�I*0<����w}�X~�� ��u���vDXU
����v���en��c��X�v�� �\��@b����&0�� �ф 0dH�E"�!A`� (	�R*P�M%� �\���Mf䔵�n���a��ɻx�ѹIy�1�F*9\h.��d���:ܶ���7'g�����ư���]��uX�ӵ��Aۜ���Z�k�+.�mch�kr�oGi�d�6��g��2]��lJ`�g=X�!��s	�E����형�^8�E��}�����������(͗f-��'���P�R:W�Y�r�(ݥe�f�-\K�%�@m��)e���@���;]2c�^z)�aC���{mv�pbݜ�@[���n��d�r�,�`��x�ۨ@wH��EH\9��3v��۬/3m�l�?���n%Hr*@wd� ��ŉ�JKP�"*0��ŀw�g�B_�9�����j��c�<(��]��V����?}7^ݝZ�<�{����x�M�Y$�ȆK*@{�K@}S����ʐ8� W�f�E�R�T-V����0�ǵ[v����7<����5�틷6���*�v0�H�T��F́��`c�k�>��svp���A�䂶֜�x�wqe[
"��\P�$�	w����`ns�6<���js����V����>��5B�z�ٰ1��`7�e�J�'+�X�d�������� ��j��I�{����}0���j7%h�9�n*@z8��Z���?��v�x�ۢ4�v��� 2��l���g���[uYc&�.
��,��;�5ۯ=�fn�'ʐ� <�K��a�9��o���5-v�������X��ـ~g�ۀ}��,�M�{��o��䤈�v����>g�ۇ8���� " V�"�"H+JԥQ	GЖ�㭭,׶�� �H�T1�m��f�>���m� ���,q�{}0��'��I
K]f���� >���^���@rj�veu�pn�㐎��#�y�ct���co��yw�u�m�ev���]��e��n*@u�1 yɿW�:}��~��d�r�+�`>�fy;�}��o�����b6�7n�7+n�.�u yɨ�`��ܟ*@�z���X��Z�ynہ����~߼Xw֬:�X|��5R�Ձ��e�ԶJ��;e0��ŀy'�����޸�ۦ�6�(��-Nѹ�]��v:ܞ�ت�[�5�^6�yZ}�U9�4��y\ˎ��������{�\ ���G�@w8�сs3E����w���=�j�����*@7>T�M��q6o=�~��$�����}��@w8� >�P�����3Vk����q'��~X�}���p<��ws���o�R�r�e��XN7��'����,�;V�AE�"*'�Q"E�=tz�:��mf���'���۲�p۶n״��4��ÜmGn�:m�wWH8���]�p�<��
s�vҦ�+� ]�݂�H�ۮM�!1�,,�oC^ydql��һ�Aq�F�Ƹ9R�z���%9�t!����_:q�����q�&��:�7g�8ݺ�Ʊ<�X6�5�Y݊��m�5�ֻ.��1��8wU��."�ظ^*ݗ���������`��'aݦL��O�յ����cW�qmr��qg��k�jK�!���Y�]5��=�rS��9�������*@zܘ���R�P���^Dݖ�w�L�\���R���`d�� �q��IDə�uWh�V^f�Fn�o������;��`���P�l��Ȇ����9�q��w���X̦Xz�%���Ł���I1J���$�`�������6[�ݲ�fiy�uw�&pPG/Z�lp��]p��ìu:s�t��^�����8y.q>H'r7I$)%n9o�;�t�>�L��u�">�1��[9�c+�������"K�Iqp\J&�j����;�u`u�2�(S&�~����r�\V�`�޸�{5��H9�@{��F���{enQD�UV�S8�Ձ��Ձ�:e��o{�\���b���"j�ݷ �z�X�������XsXcOF��=`���;G%�ˣM��X�V3b��Û��n'*��u}��v,�N��n�x�o� }&�nj�����l�c�*��� ;���s��w}p�}� �ݺg��g}�?I1J�*��g�U`�Ձה�)5"@�D(�DB�s����[��pR���!I+d��{�>�}�`{�� w�ہ��\�{��{ux�S���	�UE��t��D�ݯ�{V^S,������@�7`���V��\n���6�3�k��p@�-�p͒�%���C��ځwFn^�V�����Pnj�� =%� �wfYkj��Z��n w�۟З�.p~��`g�^,:�Xu�+�B�]V!T�m�>��0۷L<�7������>��`:J�R������ޖ �v�3XW�"4�@�+]8� s�Ѩ��TMR�$���[L �۷ ��^�n﫠?o�X��`vrbq�JyUZ��Z�t��i���N��Ѫ���.�F�a�����`�.Ga��F������?�����j�}t��@y�V�b��S�qr�������:�ڿ/(�?W� ��\ ��n%�&�n��,����`nmi`���(�5��5�{��Ylr
�c�Wm0?��o{�\ ����v�<�soK���YJj��[�r����������@N}��RH/QC��X�j��>�RuЁɒ?@f����S`�U2�AM��s���hB�*��x D
i����!h�!�,X0>��}��Ǝ c L�hDb�t��!D"E��>G1@��y#�b�H$¨UH�c �� ,& �X A��j��!1�����8!�`px�z3Yk�VGE��0�A�(�S]�Ç�;S�ë�Џ�0C(���M�gP�R0�?,!�#9ė�HH�I�'�r��E�%��j8$�%(H-�i��  i�p[K֒l��[TR��eZ�,`�u-����[Wr�Ȋ��P
���p�<�tQ&VN�pn3q�÷=�{#�2�'X�an(�d<�ͳGm77�y�n��Ri�Eƴ:���B��	�uGM���l��0*�\\�\`�Л�ڮ;6��%�֙�K0�kI�#N��J�:�;\�`���*�k�eXy6ˎD{�v�{V��s�]8���v�g�m���=��v��[�'ѝ��8�'�� �c+nM۲�#r�t�V]�॥ �퉪�y^���y���	-$7l�8鑶��.G�$�*�cN���,Sj��^Z���;UT�:�m@�GU �驴�wW66:=���@��UN�3���m�����Cn��.���v=A%�B1�{�ZR�sc�2��#�7$sc�ө���W���;j��R�Dc/�$^��M��K'[6��(�,ӥslƬ�H)�ۄ������Hf@��a6ll��I��L�ɞ6*6s���:͇^ȆW9��r�`�cmfv�(9p�S�v�K�ir��*�j�7c�m�A�S]:��ڗF����< 	MJ�]���X'�����m/�غ��Ħy�G:�h���SB(�����\�<�m�[���\�q�R����a둭��m��3��9w���nԒ���B�HOSm�⺯;-�`ѻ{z'Q�UR�ԫJ��S��H��n2�*��\�;*NM�t��!*�b�`��i]%����[% �nn���l��񐄭�8rH��:���U���Fegv���3�������*ԥ��r��i��쁩q�+��̱�g��zg�y�WL��bK�D8զyY]��
��Z�M�*�R�d���$jT6���ȪҭU]�U�Ŵ/PXֆ�6Z�i2�:�y�'mm2���i�q�L<�ɗ�������;l�nkՎ�Y� sv�f�_{��������~Qʪ��:�E#������9Pv#�6���� |�6�ȁ~D�+���rd��-�$�m�s\������=�Qg6;	+N�c�[rvƴͰsW�r9,#γW�7'n�z�-#�	�i��]s��w��1�g�'4N��(�l���	���:ŧjS�.ܜpn�t$��qz�[u��}��MlG0������*Sx�����ʃ�P��e�s�g�v�]��d}t��s���Sjsۙ�������,d�Ӳ��~v~���WF�P���: 㩎���p7���=���N|Z���k���_�Yq���Lvށ��ذ�n�߷o���}p��O�t�����~� �M@���*@z�YW�73/6��wD �M@�G ;��0���ɊT�r�mn[p?��׵`f��`g]2�be��X1�w�G�J�r�����;��0�n� �{� �Iqn�kk�$Pm�g[=����#�v�g�X�ry�۶�����>n��*�P��Gl���_߷n }�ۀ}��X{��Ylr
�c�W��jI9�{�l��H��A���]̸��ŀw�g�g������Z�\U*J�� �{V^;Vze�֖ ��\��ٖ���"�M�n�}��� #�~�5 F�=c�r��5:�
�V�m� k�}�v� ��n��q`~�h�9E,-B,*��nt9������BuX�h��%���<�<v��wYk�9,���$-��8��޹���g8X��ﳤ�Kı9��f��O�b%�b{���i7ı,N������1���s�ی�:Mı,K���t��bX�'��l�n%�bX����Kı/��gI�6%�bu�a}�L����n3�1q��7ı,Ow�٤�Kı;�k�I��;�~J �0����MD�����n%�bX��{�_�&q3��^�^$!�K(IX��d�n%�g�������Kı/����&�X�%�y��:Mı,K��i7ı,N�ž��m��������s4��bX�%�=��7ı,�w��n%�bX��}�I��%�bw�צ�q,K���\K��9��})���p�n��@�i���زsnu&��u���l��^x���w�{��Y�/=�gI��%�b{���&�X�%��{^�]ı,K���t��bX���������+�m�s����&qX��}�I��%�bw�צ�q,Kľ罝&�X�%�y��:M�������]����[�aX��ʳ����+��k��n%�bX������K�q/{�t��bX�'�{��&�&q3��_M��&�d�Wa!m3��Kı/��gI��%�b^{�Γq,K��{�Mı,�b?��'����=���4��bX�'������Y����j�������ou���7ı,Ow�٤�Kı;�k�I��%�b_s�Γq,K��=�{���������m=m.�a��.Iζ�ۧ��ٻ%�;����f`�70ߝ������qpc7͘��t�D�,K����I��%�bw�צ�q,Kľ罝&�X�%�y��:Mı,K�;=���6Pr�ZKi�_�&q3��[�g���/��01Ŀ���t��bX�%�~Γq,K��{�M&�X�%���7�ŭ�
��]��/�8��ľ罝&�X�%�y�{:Mİı=���I��%�bs�צ�q,K�_w��z�Z�Z�L����q3��N%�=��7ı,N{���n%�bX����K�FĽ罝&�X�q3���Yd���V�Sv[�_�&q8�'��zi7ı,Ns���n%�bX������Kı/9�gI��%�bAj�z� �O`�0\�.�C'�v[�x��G6w/��C�.3n'�1���V8��q�tl]����4U��]�v��.+����-vʝ��ۘwm�n��UK)���M*�t	�V��'õi�^���5� �8y�X��z�|����1D���cs��q���ֳt���)�N�MI�;m6�����V�Hz��݋۷n��È�K&�9l�$r������W�������/;�����˶�gm�V���h}=�[u���;7��v�ȝvu�۵���CB,��'���<X�%�����n%�bX������Kı/9�gA��},K����q~8���&q{o��"|�J[!ft��bX�%�=��7�D�K���gI��%�b~���i7ı,Ns�ޓpD�,K�����K�\g9�sn3��7ı,K�{��n%�bX��u��K,[�����H��=��I�8��Ų�ی��� >���^�Mı,K�����Kı/��gI��%�b^{�Γq,�g8�է���-�)Z��i�_�'ı;�{zMı,K /y�gI��%�b^{�Γq,K��{�M&��oq�����~���:6�ɒ+�zvt�M3BBS�&��÷c�۵�a#m痫���������3��Kı/��gI��%�b^{�Γq,K��{�M�R'�1ı=�߷��Kı9���O��3L�rf�g9Γq,Kļ�}�&�Q0ș�b{=צ�q,K�����&�X�%�}�{:M�lK8���wߩlab�
�ݷ8�L�q,Ow���n%�bX�罳I��%�b_s�Γq,Kļ�}�&�X��g��&��Zʭ��8�L����i7ı,K�{��n%�bX��ﳤ�Kı=���I��)�L���\^�屹)l��g㉜V%�}�{:Mı,K���t��bX�'=�zi7ı,N��٤�K�L�k�Y��,�BR����c�������k��;���;g��g=l[qvv�����#t݌��9�s�q��i�Kı/{�t��bX�'=�zi7ı,N��٤�Kı/y�gI��%�bu�[��g�1�ً��I��%�bs�צ�p�"�q,Ow��Mı�a���}�߳��Kı/{�t���Fb&"S�ux�������Kk�����g8�Ow��M&�X�%�{�{:Mı��A' ?p�|r&�\k���n%�bX�s��4��bX�'{���qp�3��1���i7İlK�{��n%�bX��ﳤ�Kı9���I��%��Rb'����q,K��}n����4�g&ifs��7ı,K�w��n%�bX��u��Kı;�{f�q,KĽ罝&�X�%�������1�i�.�LY.uv�s�.=@�����Ŷ�d�tl,�uF����瀫�w��,K��4��bX�'y�l�n%�bX������Kı/=�gI���g8���5���Uh(������,K���i7�q,K����&�X�%�{�߳��Kı9���I���&"b%������q��g8��2i7ı,K����&�X�%�y��:Mı,K��4��bX�'{��_�&q3��]����Z�v9m�ی�:Mı,Bļ�}�&�X�%��w^�Mı,K���4��bX�{��";Sr&���Γq,K���q�~��9+R�G-�/�8���.�s�I��%�a� {���i>�bX�%�~Γq,Kļ�}�&�X�%���������;(�W\Y�
5ma��wI� 7g/o{D��wX��S��������6�9�Mı,K���4��bX�%�=��7ı,K�w�Щ��%�bs�צ�q,K���K|o9�Ì�����s4��bX�%�=��7ı,Nc��4��bX�'=�zi7ı,N����n'�Ab."b%����#�J��ER�RUU\/�RB���=���X�%��w^�Mı�0�LD�k��n%�bX����:Mı,K�wߕ��i؊
!�fq~8��Ēg=�zi7ı,N����n%�bX������K���LD�{�4��bS��]���_Ʌ���Q;m3����+��=�M&�X�%�������Kı9�w��n%�bX��u��K!I
H^���yO�z{s�*�U
h�*�"�܋rb����0��q�C4c�v|]�z�2iwh�E�H�M�Ae��s�=X�K	���a�rOj��Lb2i�cv�������)�1��V�:�ϊ!�khF�7\J�	(չ�lupc�ϔ8�nn�ҩv�C��LP �lg��e5ųl�V�<����&^��`5��c��2���@b�s)6��:y�U1�M}p`�8�3�8�nq��.W��=�흊�z�`���6��X���N��]s)B�D���d-��|q3��L�����n%�bX�ǻ�i7ı,N{���+��%�bw�צ�q,K��ۿ\�8I���ߛ�oq���w��n%�bX��u��Kı;�k�I��%�b^��ΓqlK�w�������9����ߛ�oq��N{���n%�bX����Kĳ�{��gI�Kı;����&�X��g�Ox�����*�nZg㉜,K���4��bX�%�=��7ı,Nc��4��bX*؜�u��C{��7��������G͢�*�{�7�ı,K�{��n%�bX�ǻ�i7ı,N{���n%�bX����Fq3��]Ӂ����K,�v�N��k'gn�۸���q�㧹w��vb�_����}�-V�r�Ze��㉜L�gg��8�ı,N{���n%�bX�����&"X�%�~Γq,K����򶰭�AD7l�/�8����u��6U�
J'h"0���m>���'�ֽ4��bX�%���7ı,Nc��4���1��'��Y3�2g2.s��Mı,K����I��%�b^��Γq,��=�cI��%�bs���&�X�%��n��d$��i�_�&q3��W�����Kı9�w��n%�bX��}�I��%�bw�צ�q,K��П��v�krۜ_�&q3��9�w��n%�bX~P���|i>�bX�'��_��q,KĽ罝&�X�q3��v)�(�,E*�mn�ѭ�,m��	D�D��c��y�ۣ����x��|�8�;d�g㉜L�g}�����%�bw�צ�q,K��9�cI��%�bs����Kı:p�ޘ�qss.$3q%�M&�X�%���^�M��C1��;��4��bX�'q���i7ı,N{�٤�Kı=�ҿ/��9)]�Wm3����&q3�g}��Kı9�{��n%��1mS&�&6yD�B��>�t���
D��D0�@	�c�G���9Y`	��`|	�!zjJ	�
��B 8f��Q����# E&��ā!�Q��_�L�Hj;�1�
`;����LJM"Uke*:ځO�q��-����`�
Ty� ���|;0�O�w�d��:��U4�TK�Δ�� aC���D�Ms_l�n%�bX����Kı9��tOg&qc���s�&�X�~"w?�~Ɠq,K���~٤�Kı;�k�I��%�bw���_�&q3��_w}�Uju�b(@�Mı,K��i7ı,?# ��o��}ı,Oc��cI��%�gg��_�&q3��OV�~���� m�ɰ��@7v�ݫ^w.�����62Ç	�V�q9]e�4[Vמ)��w���oq���4��bX�'q�{Mı,K����	��%�bs���&�X�#8�ۮx��X�,j�[L��q3��V'q�{Mı,K����&�X�%��w�4��bX�'{�zi7�,S8��B�#��v�h�8�L�g����&�X�%��w�4��bX�'{�zi7ı,N��4��bX�qj����X㶊X�Y�_�&q1!bs���&�X�%���^�Mı,K�罍&�X�_��*"���8�Nf%����7ı,���/��Y *�;Vq~8���'���4��bX�'q�{Mı,K���t��bX�'=�l�n%�bS���K�-懿�NO�B�#�ЯE%��ø��Eڬl���{:��-,�����'�-�rR�d��g�8���/M����q,Kľ���&�X�%��w�4��bX�'��zi7ı,Ns��Og8������q��Kı/��gI� ؖ%��w�4��bX�'��zi7ı,N��4��bX�'��g3,�3�4�K.3�&�X�%��w�4��bX�'��zi7��,N��4��bX�%�}��7ı,O�;�,�͙2e�s�d�n%�bX����Kı;�{��n%�bX������K�T,N{�٤�Kĳ���qz!B�IcVB�g㉜L�q/y�gI��%�a�D#����:O�X�%�����I��%�b{�צ�q)��&q$�sE�����mT��n�K�B��<��=�ۏ�R��p�j�%f�d�у	�m�Wn+�n9/U�^n���bm�8^��ru:Q��K��|n
wF��]�a�����b퉤7d��u������U����n�
��\5����nګg�xڻE\y�Uv�c�Wkq��O[��St[��ޠ�8�8�iv�����6漜���xzѓk���{���{|����X��'$��<z��Z�:]v��f7#aۣ�j��]�;���Mۧ&;d����N&q3��O����8�	bX�'=�l�n%�bX����Kı/y�gI��%�bt�[��g9�1�\ۜg:Mı,K��i7ı,Ow���~~���%�}�߳��Kı/�~��&�~@"����bx�'���󋛛���s�I��%�b~��~�Mı,K���t��c������~Γq,K���~٤�K=���������H��R�[�w��,Ľ罝&�X�%�}�{:Mı,K��i7ı,Ow���l�g8�����=l rESL����%�bX������Kı@{�٤�Kı=�k�I��%�b^���q~8���&qw�����mU�Ka"l�F-s���s���񗇎D�aN-��Ol��҅b�����g8���o�i7ı,Ow���n%�bX������Ϣb%�b_���:Mı,K���S�fndɓ.��3I��%�b{�צ�p�l�q0�h �bb%�{�}�&�X�%�y�{:Mı,K��4��bX�'��b��W81�f���f�q,KĽ罝&�X�%�}�{:MıQ,K��4��bX�'��zi7ı,N{��-�7s�bY�g8��s�&�X�%�}�{:Mı,K��4��bX�'��zi7İ�;�{��n%�bX�;��x����sg6�Γq,K�绯M&�X�%���^�Mı,K�罍&�X�%�}�{:Mı,K�	�SS�s���a�Xd.y��n�&8.���+3�9�wn�N�ۋ��:펳I��l6�����K��}�M&�X�%��s�Ɠq,Kľ｝
�%�bX��u��C{��7����8?{��jd������,K�罍&�X�%�}�{:Mı,K��4��bX�'��zi7lK��;.��sa��$�K��Mı,K���t��bX�'=�zi7ǚ�&D�Oo���n%�bX�����|B�����{�)I\Eˌ�I��%�'��zi7ı,Ow���n%�bX��=�i7İ?���z��)!I
HY��%yISAK&\�s���Kı=�k�I��%�b{����Kı/��gI��%�b{�צ�q,K��(!�z�~�.��ḋ��=�z�����onwE�y[��N^rA���&��Qe�_���)%t����bX�'��1��Kı/��gI��%�b{�צ�q,K��}�Mq~8���&qwu7���A�[+��Mı,K���t��X�%���^�Mı,K���4��bX�%�=��7����'�y����\\�0�qsnq��7ı,O���M&�X�%���^�Mıľ罝&�X�%�}�{:Mı,K�$��o9���$��e�s4��bX�'��zi7ı,K�{��n%�bX������K�����T�<����k��K7������8?���|Z�"n������bX�罽&�X�%�������Kı=���I��%�b{���&�Y�7����������W=��NJ�y�v�]՘��9؎<V�焳Hb�^5���=�9)��:Mı,K���t��bX�'��zi7ı,O{�٠�>���%����oI��%�bs���&33�.pLɉ,�3�&�X�%���^�Mı,K���i7ı,Os�ޓq,Kľ罝&�A% 1�8~�)��bL)��e5�O���A$N���5�?D��}�&�X�%���^�Mı,K�=�Od���1s�38ɤ�Kı=��zMı,K���t��bX�'��zi7İR��wߖq~8���&qwwĐ$��u�-�.3��Kı/��gI��%�b{�צ�q,K��=�Mı,K�﷤�Kı5����`�I��9�y[�J[X��N�%u���7!ݞJ�ڋm����뇨D�vtדu�vT�T�E���'�Y
R\v��[j\I+�/�,���;R�m`	�r�$�woWk����7`z���l����q�\�9�n7R�ݓ1$[�l	�c�'k�9@m����+`7��:�hꄀ\��q�
h6zQY�Gh\&,p���4tD�
ڛ&$�s�Ɂb�nP�uۧ��u�]����ݛ�uXx�=]v1��N�N���{�_Α*ܑ$������d�>���Kı=�{f�q,Kľ�}�&�X�%�}�{:Mı,K�I���sssq!��ˌ�i7ı,O{�٤�Kı/��gI��%�b_{�Γq,K��{�M&�%�bX���[�y��nq��ss��Mı,K���t��bX�%����7���LD��k��n%�bX��~��I��%�bs��=�fbF��-��s��K��$P�L~���t��bX�'�{_��q,K����M&�X�%�}�z�㉜L�g��~V�D�@d�s��Kı=���I��%�b{���&�X�%�}�{:Mı,K����/�8���-��$P�$���Q;.��^��{m�i�mck=ˮ�t��.JH0}��_�;�4Z�덦����{��7���{^�Mı,K���t��bX�%����7ı,Ow���n%�bX�=�J{&)��9qs3��&�X�%�}�{:M��H@jbf%�}�o:Mı,K��4��bX�'��l�ߛ�oq���?���)���Zi���n%�bX��ﳤ�Kı=���I��?��������&�X�%�w���/�8���-[�~�v�G]�\�I��%��R�������Kı?w߶i7ı,K�{��n%�bX��ﳤ�Kı9ä�o9���!��ˌ�i7ı,Os�٤�Kİ��E1���gI�Kı/���t��bX�'��zi7ı,N�L����� $&�2v���KI�����9�:^�oNn�w\kk��wG�#�b��&�X�%�}�{:Mı,K���t��bX�'��zi7ı,Os���n%�bX��=n{��d�g9Γq,Kľ�}�&⨖%�b{�צ�q,K��;�M&�X�%���z�㉜L�g��~VWcb(BY��:Mı,K��4��bX�'��zi7�+�W@�@�B*�Qi�쪹�E�f8A%��P��?#��!�@N ~� &�_����n%�bX�����7ħ8��~my2�[Tm�q~8��g� b'�߷�i7ı,K���gI��%�b_{�Γq,K��{�M&�X�%���ԧ�c8pb�..fs���Kı/��gI��%�a�P(���߳��%�bX���~�Mı,K���4��bX�$Zrr[�b=r���H�v�u�ۦޜ��N5t��\)�Iqכ�ѵneÕ�]��_����7�ı/��gI��%�b{�צ�q,K����M ��bX�%�=��6q3��L�ջ��б�m��ݷ8�D�,K��4��bX�'��zi7ı,K�{��n%�bX�����������8�W���?B�]�v�J�7ı,O߿k��n%�bX������K,K���t��bX�'��l�n%�bX���[�y����9͹��f�q,K��9�cI��%�b_{�Γq,K��{�Mı,	�m���G��`f�A�O߿k��n%�bX���ۃ��cpL��3���Kı/��gI��%�bs���&�X�%��{^�Mı,K�Ͻt���oq�߿�c��߭l��t&,�����tBY���&ܹ��1��s�,�v�sl�0\ɉ,�3�&�X�%��w�4��bX�'��zi7ı,N�>�� �%�bX������Kı>ǯ��]-#����8�L�g8��g��q,K��3�]&�X�%�}�{:Mı,K��4��-�bX�=�Jc�9Â�����s4��bX�'y�z�7ı,K�{��n%�bX��u��Kı=�k�I��%�bs���9_q2��w���o�w;ݏ߿~Γq,K���k��n%�bX�����K�[�Ͻt��bX�qj����X㶊X�nۜ_�&q3���w^�Mı,K���4��bX�'y�z�7ı,K�{��n%�bX�8#�N�8>HN|����@���7�JȋEpWS
F�Y( �@
�a Cf(o��T��&YTH�R�3�2��$�B0P��!�>��Ld $�!���Rp�3)�&�@��c[�CL���D���Q�8X+ß(�M|Ǫ&����!�%¤�����Ċ�-�کÀ���A!"�m�  p%�niz�mm �BA���m�m�e�Md��Z��X�/1�T����Ϋ����tCYg3�vK�K�E���\Z1�ޑ!:��<��-=�� !r����FVͽJۂ5�g�5mF:UlֶmK̎�@�,�OnѮ�;<>h1ElmN��1��bjlnx^:��m��r�M�U�ts3��Au\bǝ8^�N���;N9:�F��Z���<�up39�mz�KNr#l��������M�j�-���iP��+��)]#J�Q��j�s�y�X*�����:71�vl�U���"-�.��͆� m�V� �]�J�X��m�l�SV�r�\d�-͍��ѵ�$�m�6Z��N7\�lxY	�.{WF��ԍ�C*�� �Z�Z�wY�UJ�r�8VV�L����N��8a�R��	���!<m=bEi�-#��s�՟SX��nU�:닭�RxW]��Xظ��ef2�>��p�g�l�ݲ[ؔx����� #�	��y�u�i����#qvp��a�^�:u&s�H<�;C1lr�"ݯWnz�j���e(p�`��v��$��s1fQ��K,�/B��q#�������t��[wk(����* ����U�X
q�_>8+�]�;A�P�E͌`U.����aj2����ke$t,A\i(ɻ3�P�z��n�$Z�\qƚܻ*�ԫ�*�pW��]����I�n����(jU8z�Ōtڮ��jM�˒��zr+c�W'#�LXq+�ۉ�FRZ���b&eg]��ݭn�vL�9�d-�k�v����v�imٍ㲙 4����M���Ay����lut�ݩR=��,��:����B2۴�m�l��T��P�UWmP�*ħUCjZ
Zt@W�X�[�e�mV�Ws���lFDul�`gnàz[���KÜ�v	f� �sm�$Ř�3z��\�"+�M�T>@��4;�J�������h����D�	�*+��P�h��o�3��9�1#	�ルɻq���4��A6�`��N4N�tvz�R����+i�{����$:�bV�˴���arn���sգ�/��AqLPgrj\dd��IprKb��.���;:�<X��si%�ڋs8���p��{Qn�=&��2Y�gLZ7�:�m`Z3�L^��v���e��ț���!��X�n�i�5?�{����q��[hq9긳�'-;Z
��u��;�����۷k>�t;���/$�J쪖Q�Oq|q3��L���צ�q,K��3�]&�X�%�}�{:��蘉bX����4��b�ow���Ӄ����UU��~oq�X�'y�z�7ı,K�{��n%�bX��}�I��%�b{�צ�qRı,Nc��=�6��%3���7ı,K�{��n%�bX��u��Kı=�k�I��%�bw����q,�g8����[�E)%����q,�";���4��bX�'�ߵ�i7ı,N��4��bX)b_{޹���g8������C+��u@��s4��bX�'��zi7ı,N�=��n%�bX������Kı>����Kı?=�?}p`�q���\t�\r�^��	ؖ��&51��Ӹ�,����71���s�����9�S炼��}����oq������I��%�b_{�Γq,K���צ���&"X�'�ߵ�i7��{�������eb�q2�Q���x�,K���t�����~E >�"}����I��%�b~��zi7ı,N�=��nbX�'Nv�1�c9�1�\�s��7ı,O��zi7ı,O{���n%�bX��{��Kı/��gI��%�b}Ӥ�o+�TQ\�j��_��$)!n��p� �,K��}t��bX�%����7İlO��zi7ı,Nx�-��"���붙���g8�Żw�8�	bX�����߳��%�bX���_��q,K����M&�X�%��M���8/�+h� ����|x�u[{n.ל[�Fݧ�OV�䛠fL=6��q��n��%�b_߿~Γq,K���צ�q,K����M&�X�%���|����&q3���'ic"t��3�&�X�%��{^�Mı,K���4��bX�'����7ı,K�{�8���g8�k��+����\d�f�q,K����M&�X�%��羺Mı����� 0H�H�GL0 p�� ��D�K����n%�bX�s��4��bX�'�wR�=����nfq�I��%�E����{��Kı/��gI��%�b{�5��K����B���
HRB�u���*j��.q��9��n%�bX������Kı>��zi7ı,O{�٤ܶu��`{����孖"�����Z� X�#^EꂨΔ�Ӄh���ط.�^N/�"�:۶��y_��,�����./�{޸ڵ�[��R�:�,۵`d�>XmՀ��2�&j֛��I-�'K*�<�}0wv��J�����ݵ`vz�'4HEp)J���6�X�S,۵`�X�\�+�~�� ���N�d"t���t��I #�- I&������]�@��܁]ۛv�^ۇ����ێ�Wq&I�f�zYiUmڰs�m�����K��F������WK*�7����q����}�+� ��ŞK�Cvy���؎MM*�U��{��X<T�=	L��X�����=�X㶊X�nڰ��j��7wmX��6�Q��{��X�Q躢yU<��r��TX�j��I�z|��V�T�T$��&���r.]Z���[[ta]n����%��7��X�^�mڵgD�\��ݙ�bǮ�q�[n7='cZ�z˞y�gt4A�A�,i��iq�욲+���9'1c��kk�m�v`�n;l��tW5�,rkۗYy��R���p',���N;bw��=gs٣��ț�'mZ�v���Ïu��k(61��Zΰ��ۚkl�\��Z�8v!��x�v^�����z�s��}�U��d{n�fݒ"}� 2O�U����v�6CsR�F�i��������������p�T���ݭ,�rOʩ�+�JQ�� �M@zJ� $�o`����N���:%���t�7v釸����{� �;��]-��n�耒l�� �MA����<`^�5�E��t��{ۥ�6�XͧVn�`~K82D=b�ԜOD���t��0z�\�E������ ����`�.`zu8�tS��n�Հ|�u`6�I} ��֛O�\��Km�p��ۇ��s�)$�e��� m��3�!��nR�R���wn�{ۦ�g��\ ��^�ں�z��NKm��wDx�	$��*jI�@s��qkU��MS 7wn��'����z��;��0��0��mU�u�� ��'k���[]�+w���yq��)���[%h��**��Y�hd���յ$� {$��v92��oJ��)�U*��L�D%	%������M�{��XͧVO(���rI���*��39�l���+���HP�O�PID�Ң���|�p��� ����Z�m�U�mv��Jgwv���j�m�,�cx� ��Km�p��ۀI6m�@I���2���ݬǭ�fֲ�W;�g�d���6�3�s��ݶ+*�L�=��{����o�^�����#u~ln�i`d�>XmՀ|�u`u��3�-$R�\N�� ���3��s����zP��� �gK���g��ŭV�L�l/sq I��P���	&� ����?}���u�Țu��%�qB��{W����^,���D.�DDO��͸Y��CN�["|��pݦX9�� �u`|�v�%
F6�0����v���aïA����-[��b��qrkB�8��G������sߕ�{����QSEU���� x�X6���`uu�S���S�»f own�iڰ:e����z�"�:ӕ;|r[Ev;-�>���`ݺ`�� ����F�-��RJ:�X�L�39�l�:��J!OwV����^�夊Wk���`wf oqՁ���X�ڰ>���92���K�����g���/�ꣶ�A�d���Tp7��u��m��x��nq!��H�7&�hp�J��m��c>��#���9�v{6jIr6N�U�������gd��&2�������-��Q)��b�È�������ݙ{]�pu+k���+�]�aT��v�q"c�)��f�O��W��ƛL;f�n�;&i�]n*���Qy:�r�n�q��w��{�[�|8j�#�9��=���%6�/a�my��Cb�.tT��u�*��R2�vY������`>�k�
�A�=��{jyx���41�p�ո��w��v`��s���gY����]VF�ir����j���|�aDz����X��_ذ_wq�S���WK*�:���9�@zJ���T��d��w�2R�U¦�� ���DG��Y�/ut���,��ـ��΄�*V���+���w����ŗٻ-ԯoW�3�=����9`��(�c����� ߻����f o�ۀuu˴r�,��L�jI߹��eD	 ��,8&�a���&ﹼh��\�t�g�8�g|�פyi"���t��^� o�ۇ��o�� �wذ��d��_q�����s�J��>�?��@NqR�9�s�^�5]q:F�;n��.���� ���0{�p彯�Ȝ~����,1�ۦ��N/'��oa����.���%Řl�ww&�b�ۮ��dMIIO�����,�q�@�j�͂�H�+k7J�/w�ޛ�H<r�����u�@>q,��\l7�Y�9l#u:�����w�ԓ|��L�]���2!��3���!�䃃F�lJ�G�k�
�cĀ�S HH�% �c��WY(�bk��"\Mc&��������%�=% H�ӱ�$T��݆���D�)�v�� ~��@*�>U0�ӿg�5$�q��I7í=��$��:�ۀ~�V��;�w����=�����������
fi{Y��|��9h��@y��������m���� $&�1R)�T�ꕦzۥY-�}��{��w<���F�!K\N�U��o� ~���?w�qy.$�����,^��Ό#*t�m z9�7QR�x�=��ei���4:���n,�wqa�q7���������V��t��8�r�U+D%������ٰ�:�5"u(@�ߕ��n��R�P�$�EM�V��s`y(������Ձ��k ��{ �6�mTv�ܵ_��w�m�=�����j�qFG�N����Ѣ8W\��ӛ��ͣ2�6��j��T�������?uu�����G]�[p��v��Q�B�p��Z�3y�� }�V�˴r�T���V�v�~��?�g���۫ذ[�ds+���r�U��S�Of�7Ձ�bv��n���C]
Ȫt�� ߻� �
[[���ZXg1́�Ga ! A�
*�X�q��Z�d:UL!�c�&1$1��6��n%�9^%����Eg\f�O$c����lP5��L.�m��O��_`�ː���Z�b��m���V6P��J�. �f���	�� ���R��)�V#4����&M7VǠ��Isms�m�KE��hmu:#.���:�6�MԎ��p�A�
�ZQ�5մ�ݻu�Xv2p[R�ų$N]U��ewN�ɱq�g��""~ ݄ì\Bo9�ZC�3Ő�]���exv��']������n�g�Y�ծX奕���'H��-��yn+�)���s�(�H�j��4թ�]+��E-V�~�� ���x�wn��[� ���8�������m,����q՛�z��V�,Wۮ�-�n�*$vW��q�w}p��T���7�@yӺ���L�ʎMMryUVىڰ<�B�[����|`�ݸ��ݙ]��R�8ڵŝ���gN�=��9��.ݴs�٭�N��|Ԓ�[d�ƥX�ۦ���`�ݿ���W�`^��erB����f���3٬���d9A!	(��ڰ;�m��)�d�p�4J
9%M�,�Xf'j�B�K���|`n��u�[
��$�UXj�	%�f��X{^,�)��wn�4թ�]+��NKU��� <�� NsP�����LՆq7g�8��Ѹv-�E�`"�;�Nに�a/�a�
���{�M���nx+�Er��u���qՀ}��y%����, ���d�F�r�F�0~���BS!��Ձ��Ձ�e2�	$�N��?av�J�rۀn�\~��S���_�v���h��P?%�}����0����>�yv�)Uv�K�������7�@����j պ��)a)K �%X���z)�{_��ڰqڰ=w<'�;��vglv(5[Lmǐ6w��v̋Ύѷi�ۓ��ض-ml�:\�:8�M~m���}�7QRs� =����wU��)e����Y��M����o�_�ٟ͝f��M�b����[�����@>{�s���]n犗*�qMTT�UE��/BQ�{���~���jI���H 鈡U  E6�E"38J��8+ħ9'�3� |��u�,q�9Q�������ߗ�n:����2Ϳ�������I��s��6hָ���M�5�ʛ�6��綗�c���������������3w<?�� '=��� 5�ݘ�7�l���V����`�uR�� %��B*@���f�G]��J��ۦ�gu���./䒓��b�=��ŀ|ϻ	j�:�+[y����R�.8�wo�+j�\V(�c�`��q`^Q�}��5�x�>����B	B@HHH��;�;w����9�V��W"�/3�oN��t�����Bղ���O&qa�����۱��A�ܻ�:�o�#�GkU�C���pK�����_�m��w9�yc`A���隄��W&��m�z�=���/�˻��u�1n�]��R���fK'"KRM�q��q�]&��s�)bOW�f@���^�+-��+ϳ.�	�&��e�������{�]�w����դ�!��#ȗ[�5o[��0g���֌\�8x
�8}մ�NG��Ɇ��<�ڻ���}��R�� =q�@{� t��R1�*�eX���\l��}0���`��� 5}��nX�*r�F�D�9�s"�� <��掏r���T���`�鸰��ŀ~�n��O����;�ܳЕ�YZ�ݳ�@>qR���� =̘����ȣ�i�*9+�#���'��&ݘ�.�pmog��� ��%B����d�7.���@y������W���a��b�:��$<�|u�WG)�~{ى�ʯ�<�*@>qR�� =�a���W�hc����q`��,<�M�v��n��3��H�-�M>QT�?(��ߕ��֖ �X=K����yw}�+/,M�Z�U�w��075�.*@N�R�xB�>��p�-);��R:�n�V��v��<��<���;��w��������dMpݔ*:��U���V�v�}!��+�'u?em��er;m�;�j�w�{���r�`1��"!%2f���ÅUU*�T���V����e�Q
O�Q	 � VE$ZQ(�`DL����<
ܹ��ԓ|���I'Nu7���*��t���{t��v��K�a�
=
!B\����#���U�o,���D���w 'H����`ova#v�F弩���W��[]+Xs���b��������)��\1��/L�ݬ�,��@w;���T��{ ��n�7uF�-�j�	�Z���_�	D%���M�{w�`w�.����8�P�9-jHYV����75��*@N�R ��^���w�j���U�(Q:�Ձ�s�������B3�ަ��t���嶸ݶ���q`��,~ۦ o{� ����FJ;V�NGj���ewS�W'�pݙ�W� �T#�� N<�B�[Z���`��,~ۦ oq��y%	(�=��V�S>UJj�J�4��@N����w 'Mŀ|��`�Ze#+��`��p�K�f���)���V�֖��er�Wd������X��� ߶����?3����UZ�ݤ� 'M� ��@z;��HR��0��h(	�H��05����"�2T#b�E�|H>*V/�����ĈAO���-U8@�@�ӓ���PB�@:v0� �����DdӸ�t�P�q�@ Ef��*1�P��1H�c*�'���,Hp�J5����?��;- Hp��vPH-��  ��-�8l�Qmm&Ed��fE���s��́������mۮ����m��H�l�M�`��z�ճ�*.�I��W�[��Gv[m�:��a����`ル�z��;�e�\��]h.���m�Kr��H$�@X1�ۙ�%�+˞��m9컵l��S)-uI͖�z�gb7V-�a�v�v�ks��nt����s�傷;v��ڎ�Ru��Iu�m7���.o$]��.��q5�DK��:C�=����m÷MA�G�O�[�Z�% M-��I .�$m�ñ���Н�E�Wo�I��� 6�mZ7U���U�ͦ�����jl� �7�?�Ͼ��Z���:��Xc����B��ik�i��s�6E����f����7cdeɻ�Z���ۜ�[�����*�h��F&m�_���h��Y�l�Rh[u�� �[fA#c��{f�A<j�a�,�ѳv������vNR{�^m����l��8#v܅F������Q������dw:�Aͷi-�^0m��C�D:<�C
�q3-���?��Q*E��9N�/R[zݷ,�\�T�;u�1��K6E�P�3Q�Ut�Λm���^�$k�F�r4�U�@MU#��T���ȹ��p&���ظj��6�у�A��U�s�ebt]�1��:��Nb�Pg�ګ���a�m���X��j�6�f�P'd�,dڥ]�V����5���H���)V�8���t,�F�0���{��;�Q�� $���[ee�q����umr�v[h�V��!�T&�Uj(�@��L�\ܩ��	����U��]��1��_V��[�N��v��8�L2�۶mTP�����@��^�1eV��NZ^`�)�G�m��te�%���$�����j�9e�Rp����V����^Ŕa=mٔ��sœ���j��(��r�� ��E/d��U? � �ߏ
TB h��v��S"�0d (t�>���C*��T3��(܉dU�2͸Iy�5�lk@�����\�z���t`�v��rg��[i�Au�eֿG���q��;1<�q�Y�m�Fd�[�7&m�t�q�Ga��a��8s<���vm�]fqqk$tmh��rY��u���UA;�); ׭���C��
���|��m��q/Q�<�8-�9�ugd�u���ҳ���,X�bq�t͹qm�1��&m��w�7��M�̬�������v;:�۷�}J15wgu��HZ�grg[�_wώ?�{�������OC�T�?W� y���K�`>�j�5}��r�*v�rZ`��s��I)���mX����ڽ��y(P��5�B�G9m�7m����,~��g�BIL�mi`�Ձ�O��Ts�ʥ<�R�[�`7�� y��<�$����, �/?H�N��mc��`�`yB�׻_���[	/�5�ڰ����п[PM=�p/M�vӳ�Rq7:V�����9�X�J��u�Pq�pŎ�͛xnm �������8����*��i"���׸�CHd�L�?�5g��hԓ���j@��������g���$���Z�ݤ�� $qR �M@zK���wV�X���H[V��'���������v��ڰ���<��L��t2�3i G&�'B*@G"��t�j���)�*R�Gk����޲����f�R��=^�l��l��mz�a��#ꪩ��r��}�ڰ7j�o�Dz#��\�{��A��K�-d%X��W�&�,^�X�v�fA�s�;S��[X�%X��ŀ�ۇyâ�5X=*���+��[(�	w�TvՁ�]��N�	�&
�IS¹J�R����s��U���֬�T���Hs�nm�n���[tY<��X�X��^���7^ڰ���Ǳȡ�nQ�lM��Ia\+p�ܛ�n��x��@�noR�b��t����.n���*�J���mX�`�~�q`����2K$RՀn�~�!�v��6Հ�V �[�9-��;B7%X�ݸ�����7���`ｋ ��֞�,ds���w�V�	N�7�`kݵ`7�Հ�ꈀ""��l #��U4	.Cn\�M�܍�����d%Xr*@H������ s>�f L]��\�R;UպB���R�g�=�i��׌��N�qZ�[[�G ���EH�T��9ܒl��Yp�� ����8����,��b�7{���6}ݾ*��U�X�O*��6Հ�VyD��� ׾�~�V�c%��V��-X�w:lrjs"��⼭�+q�Y"���~ۦ���޿��t�,{�� �$��^.sf�ȵB@��;Ɏp땯]�&�l�D66l�s:٭��M�mb5�{#'&��뺙����;��:���$��Dp�:������N�1v�� n����m�n�ݪ�'n{vq�<5NI.���[�&�ە�p�=�F�9�q�ڕ��gԤ����V݃�Ĵ6��лl��+���U\p�I�v4�b:j�H�nQ�'q�m��ݺ��l?����}������sߕU�)A��4�۳�^�۶+��6����62nn�F��]rņ����"�����������`<n�(�]2���D�����c#�������س�M��{�������?t�6d���֬��ͤr*@N��& '2*@uw[qQ�[��)%X��L�wy`>��XyB^P�����#��9�UJl��ͼ�@;�bs"��*@o۸����ih�4�N����oo<�f�i�ێ;]=�՚�;7On)dk\��^�m�����	̊�H�:EH�ݘ~�V��岺�Br����tj���UT9�CX���z5$�����7 �7��+`�%���� $qRܓ� �R ��]��:���V����z`�*@9"��*@y�ˋ.���M��ڻ���EH$T���HrL@|��̮�XW
�6���UR8�]�	���:ݦ �����oG�����N(��2�n��IÔ�mڰ[�`d���䣼���� 7��͸��*�����~ة �I�	̊�H��s��ɵ(
����<�`d��`>��Yq�PH�"��b��L�"P��*���}���}��F���Ӻ쭪���h��0?���t��O��Rt��䘀}��Wtnnn���y�� �Rt��䘀��q`�� �[,��,���Jy�u���[��Ls��g��ӯ�a�6T?}���|=XQI,p����{��,�wf�t�Xww j�u��]�S���`䘀�ȩ 䊐8��N��!c�T�WTv�~�q`��Xys�o���`��L�.�fH�KE]�p�+v��ڰ2[|��ITE�$���!%�P@3߻;��������*�����w�� �m��}c�`cnՁ脣!���J7f{pC]U��gx;oa��a��5��<�:��"�c���S+�L��+"�U�>��`>�ڰ1�j�o���cr�U;�#�`��� ����7{���ݘ�C�Shv�
�Br�J��ݫ�v��Q2�wy`ni���{��R[H[V��ŀd��`>�ڰ�K�ߕ�j�6�g�Wl�ڻ�ͤ�& 'B*@9"��w�^..�I,�g�VڂӒX�$`v�eְm�qq��c7lQ���F�w:'z����Kεd�S�izS���"�KU�<��vBCf%W��*�����t�g��1N%,�k�b��d��Nm96c,'k<c���[��붵�GI�b��:�kgm�ͩ-dx��T�'��w�P`��2ګ���=pm�����v3��J��t[�/"j�g��Rg9Ę�Kfs��UE2��UC:��6|�5�!�v�N���:Dۡ���h5����6����X8�)�8d,�ug����?���*@H��& =��̑�*���Y	V��ş�M�������}c�~J""�cOfg��iT*��U�{��X^��~�q`��X���I6�B*�eX��B���偹�ڰ1�j�ǎՁ��3]�2�bT$r��i���q.$��ߗ�={j��m���=�.��L�臨��%�M�t�[rlZ�^���;<"O.z�=[Z��:ک�;c"�	�Z��ݭ�5H��@�1�@u9�mn��3il�rjI��5�X��,H�:PR$�"�u��������X۵~Q�	BK�<��cmJX:��v������?}����R�� <��\F^�]nٛ{Y{���u �R�� �1��nY!eN^Wk�J���,��9�__�}��qR~���W�e�p�ݡ�ډ�\��Ǔ8�n�,V�on�c/���:ەPqQ�U#��IV߻t��1�.*@9"�_<�ɻ����{y�hrL@6�*@9"����<��q��پr�V;��#�`N���5$�{���t!m!@"�� h
-ȲF �
#��t��n_�gY�B��Y�0I�P�
2��1��a B,!|����Zd$q
�a+j)H)��0d��&R�$$�H� H��f"�
i����H��� �"HЍ�"�bD ��0��@#�	:h��ǜ(�(}�>�s_/#��N��i"ؐ,�Bb0���f0�fk$��m�^?uH�$��4�FI2[�(��ddi	#B)�D�	@��� m��Ð � `��A�/�	� �y�4��z�P� )�Po{�}u��ـn���6�lq�RWj��Q/w~Vs��`d��a�[s�+�v�V
�Z�H[V����Ĺ��}�I*@9"�X�(pݫ������M���d�;k����ݐ�"�=���e����p*E8�J�(�u:���� ���3%ڰ7kЗ��ń֜��94Yu��m�^���qR9 =�%����D(�I.p5x��&h�R�TT�I�R�=������`�0�j�;�Z*ݥV:���`�wf o[�0�j��BYDK�Q
`P���Ȃ߽��jI������L�)�r�� �=
!����5�ڰ?>���Z鱻m��刃m�dIv�s��4M{X�9/�:���ȸ�7�Q���n��,�/7P�*@G"���� ���w����;c�8�����v�н
8d�� ���`f�_�9��q����[P�(���rڰ��� ��c��ȩ9�,��+���J�\o��\t�b�7�ڰ�P��%̭��`f��>�r�3"���̽��c��ȩ�rb �m�/���J|����-��']n!e�Mƺ�F���G�:⶝�N��;^6�x�s�n:r�4���)
�k��1bq�dQU��E0�O;EU�c]gp� tvB0�3��f�u�]�֘�Q����.��m`��ը�<�����+�q��/�j}C�b�	��5��m@��#(Fn�6�),��O9��trg�8!�tv��ٵܹ�H�-��uW�.~���G"�j�+V�^�"����d�n�v���s�a�QLj���9􅬩���d�~��b�?>�� ����;���ՠ��T�J9V�ܘ���|��P�H�T�|�p�e�"��-��n���,?�.7��b�>{�L�t%�6V۬�Ǜ�t�n*@zܘ��w���@}�&��8�i�mX��� ����5ΜT�m�����������A�un;m����wku�`@tv��G�}�ǔ���*�G%nKW�>{�L ޓP��H�T���%^F�{W�&1���RI߻��/Xܪ�""��$��E�w�V�����`}�֝�;#b�Z�v[�}��ŀo{ =nL@�� ��˽76�7�ޛY�H�T���1 N�P��H�ՠ��j+�J9V��v`����i��;V�����T��W�nk�l���\���q �]��n�i1ά�=!�h��{m�i��o���ڀ�N*@F�v9h�3v����в�u� #qR��� ߷n&���ɶ9Zv4ⶬ[�V{�seTB�$D
J��B��ǖ���v���uT�K���ay�����- N�P�R{�ŀw{�8T:�uU	ex�k����{��{w֬����3��ۿ��n���4j�/h�{/n��X|77��˫�N���m��pqY���dBk�=�"�n*@wc��'I������Iye*��{�ŀ}�� ߷n�廋<�a���qV��%/6�����5� #qR�u��Z�*��W����?|�tjI9��:��������A	hmU6���~��}�;�bLg8l��YFܷ ���ŀ=���������;�{����Ge�7�K�A�nM�
�n�k�V�g���1��˴��^�hr��i�mX�ݸ�N�����?|�q`��rڅT(嬂��;��@I�uH� 䊗��o��p���T%���޸��,?����X{7� ��]i�+i�J�� ���ŀn���>�w^����Z{���ʤ���IV��� ���6 �u`}�ݫ��J("��q>pI$���̵E	�J�`��yn���#�k���U��0;�v,�[�Zɘ��׷W&-ԕ�ˬ�7B����m(�u���v�;�nvq��igJ�t���5��8��.vn09�����S�p��ۤA��wq�	��O]�Y�ω$:�Qs<��ې.�,��EM�����۟����;�Kl�x�t�/�f3��l�H�@�B��KW8���%��?A��+�XV�B|�JQN�ue��^��lB`��6����Y��Gs"�⣪�GT�9V��N����`}�ݯB_Hn�ڰ9�ry�R��9[W[���$�P�R� ;�ǟ�l�w� Kcem��6��^�+v��P��g̀=ݫ���MKNJ' �NRՀwwq`�w^ w{� ���� ����
J�,��;�s`z^����i��x�X��{��o��?�n�����3�]^�I�m�Țƹ8�u<��x�F�M�ɮ���4�:�qST95G@7��Xu�Ձ��^I%���o��w�i�T6G(Vۀo�����l�0BH#�H"�U	$��Ct�X��`�V���ݮT�唰�`������?L���`w4�V��	�iU��3ͤ�@$���� ��X�u��Z��5\� }�� �u �R�� :���2�j��p&�<��m���Y�(�[]��4<�;V�*�.�� �����!,�_�o���� �R�� �j�Lʕm9(��M;U� �wq`�w^ }�� ��[� ����څaG-d-��;�s`m՘b]��X�B�Q�����ŀ{��X��ʢp�8�v�%ʹ�M@z:��ȩ�=�Z�j�Nz��;Q]n�p�ո��b��r�I5 �pI�ow6��3�ۮ��{mɹݦ4Q�;�.ގ�7�kl;�qq$5K̍��N^YGT����$� �j��T��򴽴���`���?���w���>��b�;��X�u��Z ��5]� :۫�ڳaB�ovՀ�֖cv(��r7I%+v�s�I%��IN�W���zՁ��e�BIFGTDCP�fl̸vvE���r4�V���R�� �j��T�=Ή�����<F�6ɷ�v��^�x9n��vۉ[����n'*v\Uv��U]��S,���>x��G�P��w}j���L"p�H��!� ?n����rd��ڰ3��^2F�T�Rm�ʬv;-�>��b�;��,�wq`�ݸ�M��e%N^Yk�J�?��J[{�=�`6����k~V ���⣶�ʝ�v��wq`�$�������@w��V�JDDT����UPU� �� EW� ��� ��UW�` ���A_�
��*"�*��@��@��@b*� *T��@V*� *��E���@��A *"",��H�� *����D�`*H
�A��EF� �X
�@��B� *���", *"* * *","�H
�P
�B��"�P`* H
�X�,DX
�H
�Pb��� `*",H��H
�� b*��@� *F(���E`��"� ��P��@�"� *P� b*UP�"�QH
�E(�R�",�"�
��"�
�F(��"��"� �T�� "���UW�*�*��Z ��UPUʪ���UW� *��UAU�J�
�� U~UPU�b��L���3�
=� � �����!����|> �@ �P } � �� QZ  ^�   ��  �TDJ P(	 *��P@��T�B��QP�   @��U@$\�!  �x    ���5�]u��Ѿ���������_s�k��oCp�X�-�p F�n��Op7c�%�Ƿ9�� 7}k�ܫ�I�/����x   ( � kw��͞�}�^��z.� ���[��{��띔=���Y�ڎ�r��������F��3bY���	�.{��G�{۽2�����s��� ��@ Q@
P��
w������:3���y��^�࢝�9:��9=>���{�=��y�ݳ�o<�>�޼�^�\G��
q���lӹ�����n���� zy��]s��޼�W{�ɧ��{�� ��P ���{�L��5����۾���� v   � @ H � n�@�@A͟@�� i @�OG �  � �P� �w: 7`  ��S��}@�U (1��z}rw1�n��'���[�d=7a��������zn��8 ��89��/�ޠ_g�^�����p�=��#�w�˓K�        �5���2����2 4���ɃS�JTT�h�dщ�L�0F�=U*S&J   �F� D�*��Ҡ  �   ��4��R��m#	��d�LL���)$�d�	���<�d4G��d���S�C����&��̓���}�:��߿�P�7k���*��<DAEC����?Χ��*(#��������<�@�
j #
D�3�qQ��( �2Q���������~����cm��m��m���m��m����m�lq���ol��m��������m6�����i����m����6�}a��m��m��6�m�e����e��o4DD@�� l � �EU>�@>���,@��*��@��C"� ~���@� �� >��U�}C��@D���� >�� >��U� /�C�/�U� (@���� ����P_�?@� �_���@l�?@ ~��� �@S�P >�	�US�/� ��}�绺���ĘB�(���?�#�~�ʚCM(~��Ï	w@����cCK��ǁǙ��+�0��L��p�=��ê�5����fa0�s��y�>�>n>���n�x�{f�8[p�hr�9q�3�NV&�
s���;�)����w��&\��%Кa��8�zK0��F�$ �K1]���<�#���$��4���WP�\��������ZNK�ә١�,*�=<��NoF���c�����I���$BD��Á�;�ip�aHP��H4#bH��:��Izﴄ� ��X2̅��
�3�'Y�8s	�M0�"e���jD��9�\48�z{cS8��9���#�a^��9�0��'2i��.��!B,!R"@ą��k7Is�w��l�3'd�u�x_f�p�!aRaBV\��_w{��� Bc
0��F�0��l)�7�Ω���&���ę����A�L�<�y,�tv#1���:��>>���#�4��x��>xz�d��.�:{}�ae0!e��u/K4���v��0��ׇZ����z�7nu�\�����(sκ�z��h� p����#$��bP#ȥ"����Sd�ˆC)%�뛜l�hE�Da +�l
$R�hz����4;�BmZ���I+�fd��Ġ� bF^Ρ�6<T��8����H�!����%<��E�.$ xS�@�	p"MR�|\�ĝ���%ʡ0"�����-��K�$�:cQ�cUˆ�¦�X#����q�bh��N[0�RXs}M��wݘ��G�H�(rwli��!@�U�z �"�bE�1�@���|���P!�!+��:�FHG��׊D�:H�4 brr�d K���j��ƣ����Ԓ207��&������B�ൕ�	
%
j�q*�-s��Un)�q�������e�p�H��`�C�I\!F	BGS�e9���70$��%�°��O[�����=0�3�#�@�4�N)`l��
������̕2�\�0��2��% ^�I0�� �^$�\H͝�0�| �"D�`HX;z!�G���|���$ � ��=c��ɺ�%�{���p��������;<c;�C�]�{�:�A�p���H����zL5��+��s�sK��;;9�:η�z�nw�z&�L�H"B���al-bB$4 �-C
��w7tP9(P�� u�/���]p� �W@�
|)�Vׇ��~�
z�W91��WQ؈�4�!
�9��/Yz�D$��IH��sw�P�"��MQ8��)w���u}r_i�yL�����z�Yf�J��u)��Ny�ti��AŨ�����98��Ά���T�06$�uJ0HC�l<�@��G�u������
��.0���� �#�T���
F$J�
�"AJ.p"B:f���2Ǹ'D�`I����h驀ŉٰ�O<8��H`B�	��-��;HP���GcX�X�B)R�$R`,C"R�u;�{a��!d2��G���z�H��	I$$��ﬆ7y�!(A#
`kp�>!@�(��gX�hq���;S�pׇy�]U<������H��Z�E�ԠZ��8T�!H�RL��)��j�����k�`V73���;N�{	8�	��9�K�!��4%�M8pG*�D�n�\�U����\��r%�d��H�`S$ׄ.!
���ļ<Ԅ� �����!"D��R��HŁ��H�)B�(@%��2�T�P�e�qYR\%��HVP�M�CN v�� N��;à�@:y#;I!	 D��E�X쐬`�X��"D��=u�}�s�����M#B3;�:�{_A}띁$�z�c�8F)���B�%����i�!�u��N��a@#P�׸1� T�3N^�
�h51p)�0aq%��^�\h���,A��Q�ٮ����E�!J��.m��6gQ�\B� �d�(�1����d(@���+
���K�vn�C�߽dd�e����R6)p�3D��N�I�	C!�
L�0%8$���uDt ��u��`��7��B |�0D1X��Lrc�#��f��WIF0���IT�550���۝�	L�8�H�ї��9����N�p�1NO%\��'\9rO i�6$�HF0� �1��	獺_<4���5160�s�}���&L���{�n� B��+/�Z�2)����@�D`�8B��Hu��!�+���E!D�Jd�!���2摤`ᦛ.n�4�%0ݐ!F5ӓyx	���$F	T�"Rp��B�]$.����+A����d�C�E ��Ǿ�S4V R0CÄ�X������@��D�%XS���X	�CB0�5�S���4`A��L%0���"�1�-3��0`h�h*�k�qk��8n�����tǣ"jv�m�k����$�]� :�u.W�5��78�^���	sMcLq�B��5%0�h�s�y{�מy'����%��P��	TÑ��u�{�++� J��+���vwN��9�Jd$�a�:��a�2�(c
d�,jB��b����bF�� `������HIYp���>c�vu<	��@$ux�v�p��˧1��Ln�Cw��tq|a��(J��tۺ�� @�E����0����i���\�i�\ �=�2��1�N�i3���l����NS.��Z1����$V���1!SM!H��6HǄi��S���y	MZ� �B��zfZXR��#��(1�Q5�a��*b%X!T�`�
A�c�κ�\���U<�/�36�	H�w ]�K;e�7S��������l���v�a�i��۝%��z�Ԛ����;I���n3������u���z
��+���&�|}<�p�}=��ִ�fl�s�0�~���������!�JC��zd~��	��?+�������I$�I$� @              �            �   ��� ��l �  � @��  l  l m  ��         ��                                                                         ��,��n���$�5��m:�@�`Ѓ ���]�cv�j�S[p �%�-'6%rT���c���Fݮ-��p�v.��5�zy.��V��CK�#bw�_|� �(�U���re0�K�,Un�_m8qͣiŢݩ����?-ٻ���.m����"����F�����������[��DK�]�6Z�y�v������V�|]���0A���ڶ�tl�i ccb�8j�CL1v�X&��ӥ�r@�u���
 m�`'R/5`    ��t�j�V����p�r��Jٶ*krڪW�Ca���٤$M�S0�5T���;m�1��d��tm��A�ŉѤ6ZvN�V�b�	VRP1�V�j`m� mgJ��5k�� H׵�i9��mp ڶ���}\�a�u�=5[1�H|�}�� ��-��u�`     ��(-��� � l�	ޤ��/�ӎ  � O�����cm����pLR�[]q�kg]m��6��,��\k��$m�l[�m� l�H���s m&��]��$�m�m��|h imh�`�mm,2�` �&�[AUU@*s�L�6U��j���  ���  -� �$��kj�6H$m&� $rIe��[@I�V� ��E��` ۪���V�q�l�l��Lk��aynVU����6ٗjy�� VYWH�U��W $�m�[[lh�ڴ�h   I"�9%��qŵ �WIW kX 6��H�  ��YZO$�]���h m� �`��`��Z�u�m�� 1�n���`��m��
4�8�`���Mmņ���lm�9�R���s�k�*�Uk�t� M� 6�:H�j�e䡗aۨ 6�U�mI�i��-� ��e$m�V�������[\�^� p-6�4�*�����f�Uj���(
����y��R�]K�+T9iIn��6�h ���\�m�+�,�Qx8�f[x�k�unm���   6�+r1]UU.9eZ�G0 �kv���H-��snx.��s���Ksdˊ����m���i-Ƨt��N�v�+k��e{L�+rJ�9�P�*�]mTZ�����(�p�UD��m�p-�ӕ20 -M%6d�GrF�6Ͱ8��À   p� rT�E�����k�m��t�-����2�J�Tu���Uj�mͱ�k� ���&�[s�
Z�Y2N�y������U��=c'՛��A�pM�^�m����d�$R��n��дZ8�\��>�lXe���m�qJiK��@r� 6��kh�[�ѱum+�@m/-u�t)��m@�[USm����  � 6��% id�:F�[@ �Ƒgm�m�  h ��I� � -�8���]r�H�m���H彯����(�k�޲�n;.���I��v�aNk��p���|l���0�  l �κ�^�kgl��ː��s���\W[��brmsvh�&�h[m6   &��V����_��|M&;m� 9"�i6���$d���Hp  m�m��v(-6��U���  [E�B@I�l^�o���i� ����@l     �V�m' [B۵u�`�n �`7Z�m���Em&�  .�Y-N�鰐-� gA�Aml ��ꪔ�U2mP �[��[�Z�[�-����@-�H �� $�Z�����@t��p�ׇe�c��s[Ā�g�� �Îj[u6�p	 �,�h� H�j�WtK4�>�}� p��-6��$�:�Y�M-���Pi$�?g�|e�����viV�ڥx��̀[Rܒa -�J����yYP �gj��v��s`$  4U*�(Ԭ�UT K�-��`ۊ�m���q?T��=]U�=��-bZ��yU]��6jr�UUS��v�����t�:].m�]6 �-�ֆh�����ZV�t{n􎪪��B5������!t�l��@Ÿm]����p/���Fh����GjҜ����I��<�·=��v�\��2l��N�6�Sr�E��Vc�;cS�PM�����Nv��$�hm��$۝�7&m��$��q#�lհ	� �� ��[��y(�Welav��������@ �}��8�������n�Q�dm�(   շ��[Y @8%��Ͷm���8tQ���8�m-���8�N �,���-�^���     �Ҷ -�    	   �v�5� m� 	 �����Cm��p�`�� ��[D�m &�M�   6�6�1' 6� Kj@  8-�[V�m�   -��֐     �F�(��/[��O�}�m5�oP  �-��� [d$p�A�ËhUa&�i�  $5�h�O2;6�`  @    ��v�     m�O���8ݻp��M  -�   ��&m���a���  -�  �        �A�  ��`  k�n�u���.�i��֍�{�m���"�FJ�}]z�u��i1$�  8�8���   ����'���K�f��ӧ-�:6��.�[A�	 :�zԂCe��Srl&��&꺥vj�YPֱõ٭��[��VF�ZH�[%�!I:�L�V�6��DG��]"�p�P�  �a�m���v�@ ��$  h  �v9m�KnZ�V]�V��$�.�fm�	�� m�`  m����mB��w��>7�l�v��9�:��`�����u*���` ��n��m�e�2E�D��@� ��k4�$���ͷn� $궒�'[F�6���-lU�;+*��]UR��O-��8u��h�E*t׬���*�V^�]m�FC� p�^��`���K��`��ﭒ���`2[N X�j�  �X� �ci:MS�� ��*�$�P��ڗ�m�
�Tl.�F�5�����*�u[U�d�e]�n��[h� �p m&ܶ�   �[y"D���h@���Lp $��.��$  v�  z۶�M��9�p��S��  ��"�k,W]h !���R�<��<X��U� �d��cgC��\�T�s(�j�9�j�$�[A�m������K۷k)���-� �5[�� h6 R6+e�(�]D6Я.s��M�?7��E����� "#�yA?x~��@����=s�K!J$��HB �"!@�p �,$-����IK�Xe�� 6H����%�d���D!
@�JR�@iB����$q�!B�!B �!B�!B                        �H���HH	! '�����Q;AS�C�b��G�x/�D^�@�S�H(��Qb
�� �a����p�h(�GoJ��XAA�P��C�u�s�:@�F(��@�C�=�N	��`�Ј���@08(4=@;�A �Ly�� �w����`tb�X�Ӄ� {�T(j���U��OS�q4C�V� #�|S��҇ʛ=q�rB>j���(� J��4C�CQ�U
`�v dP��H<���p� �@�_PG�=:��� L%�2* z���)�� ����1P=*���8(��X#1ﰢ�� Qq Ꞩ���TpY�%+qS�� �p� ����}��HI$�     @                                    ?/�K�@�A?� ȁ#ۿ}�����%)�۶�	���u�R�% �5 �X
���#R*X"QP $B
�UX(�Y̙�l5���w��~]���z�1�����������O�H    $ �� -��N8$m����              �"ե&YT-�9{Wn�f��h��>���#<���ـ�Z�ԕ1�-�b�ǝ�olKԩ�tu�6����\�q��*�\h1��v�`n�%�&U��i�lmB�*�B��[A���ͩ��P&�vQmQ��MJ
Nj���F#C�J�����T�f��2�֪��Mrp)�*r�\�B*�lT��T��w���[�$qX�i�cB-�G	��dC�n��n�U@�v�E�&�Y�A��ںZ�F�D��ν��Y�+T��
�\���PkS��3�&^�Y6`��	���m��uΓ���*���N	G<O&KH!\�P��S#��7F�m����::r5c�����Ʊ�D�˳=7j��J�8m���
��Ű�E�b:����<p���V��;�u��%e[�؍������d\�W��h����p�#����FҲ���7n���/\���+m�����z��]Z�Rc�Li�����cN�����ڝuUm'dح�
��؂��:�[U!+U[ud�Gm��>g#R�"vz�mC�����m�,��	�0�5R�[-@PxfVRch��V����4�a�L�ƃ�:vxne����ۯYT�I]C�ۋ�frv����tJʘ��S�vjj�Gm�**r0�qI��Pˡ���q����c�����ې�%*2����8��T�J����H���)GV�f�]21������l曃����7swl�Ѡ����E� (	я���1D_�;A���� �=~���]�����m��X  Y׆�tP�%�k��W$�b�If�%2���7�11��8�l\�.��:�2�6�+�k[Y؍ꚜD���H�㜄v1���=rv��m�s�7�&]��-n;9��a1�g3�FS�g���Y�U�'s�v䎎�-�q����7i�<�)�{�w�^�����Ԓs�%ɘ�̤�Hr[&@G��hN�0���s��&��ER�n�f:�g�"�ޡ�p�ȑpB�<�O�qi���;�t����^��h8�O�ŧ��X;���˰[�Иj �1�.]��]!�`�T�}��t%*2�O�� �7D�>́���~i�D�6`a�D"3q��컚nNh�әM
)[OX���j�ٮ�w~�>��O'��O~� �4j�0�s�^_g����G�Ԋ<;2���}�����J�a��I�<�]��Z�@7��w%��I��*����ipv��>��;��O�l��G�#!��ou��p����wq�ݾj��"0�d�тj��9;�۷\E�\��\[�Qf-��Q̢�N�����X;��ٻ��	��3p�v�l�݃����b�^��fi"��pv�@v�]11"/%��������dD����݃����6��p]ڵ8Xo�s���}����nΑ��DRQȿ�b(�F[ې���L�ڶ"�&v����e���E� �nʞ�]����탸�<��sj��m@K��{:s���Yq����Y��Km�63T�v�C�8av�묩��ɦL��R�!$�.�]�C�u�x & �;1�1 r^�:�F�J��H�/5G/+v�B�8c`�˙�����k��&�ذ�
v��˷�u�k���\��=r\72����zs-�3�Hf}�A���,Ĝ0(�f����;�`v��4�|p8��Or�;�`f��+I�$mSQC���;���v⧟|NmQ��M�Is��݀xp�����z��>E��%Ip����FTC L�`��@t����`�q2�5S *1P(	����T��j�D���u������`  5�iW���V�[2񮍽�Xs��,�Cv0���&\N�e�+t��Fؓ\������d�fvM�R g������W,�8�[�tu��z�۵ʶ����lbڹ�]@�+�mV�;PS�b��U���M��;�6X�<�n�ȕ��{f鈍�c�W^����O����G�m]�b�x��ۇ�h$�m���3Xլ�w��������^ :�.P�IH�*RK���ܻ��f{`���\�`nv݃�[ �7`�*y����*Sp��k�DH 1y��/7{�ۜ1�ƇA��8K1��� �7`�}��w.�߭�w�fT�+a"p���*2I$�%ƥڬ��t>(U΂�j$�������#P5:>�O'�`��`�����}�n���)Q��<�f� �qX78��x�.p��ܼ��i�.t}�v3���>�Sə�f�&�ܒd0�9��_z��ə�;����i�))D%R��A�f4Ds1�v��+W���D�c�Љr" �-��!������.�W;4�]6[L��j�]ߋV��WO-݂�X�3��M��O�-�;��w%�Wz��9�J�H�JNN�f��Hz:8,J�>Ͱ��S���#Q�:.-<������}�ZL"D�$�P�胹]<��PgʞfՅXB���!�Ċ2���ɛ��h"�
��	��2cNH�s�� �݃�����3V�jI
2����~��#��w�� ���kI���%T�U�̰w���f�1��E���<��t�y��w�g���R�F�E��y�M�϶�UM��d���ק�탿*y����p�T|)$&<m��M�rly��m�����WW���g2N�.nR{�`�ʞfnA��O;�n��F�*�ܳ� `��L	M��ƇH�ևj[��"R@�qC�v�ۖn�;��Ŷɍ9"�'����-��*y��>9���jI
"c�n�>�Py��z>۰�m֞ȐB�bJI$�H ;n���]E����c��\v��is�������jJ9��`��*�t�ƀ��d�5p�jo=�u�Wks��L6�i�C�ֳ�ݲ�d�k��.�۬�̖�tt��L�1ݰp�ms�vŌ�֋��;�v�mn�W�o&�
5���B�A&)cL�\�/UT��v�u���;���������u�9n^n;D	�oVƧup:]�y�Ĝ}q��
�(a��0f-"� �� �l1��E��2��`�� �l�Sϰ}�QP$ی�K�m��`�ʞfnBp���S�F�탿*y��w,�F�10�q�*t}�O=� �oG޻ ���4���m��UN��n{uV�]l��m�<�����s�I�ܲE-�jʹn�� W�6��al�˛�L��}��C� H*B@��;�����ɗ/E�I{�B��7"��Y�1S�v�ڭ\ߴ���1C�t}�O3.A��O-����\�`n[��j�`��O=��)�0���&��r�fc�a��f2Y��� ^Ӂ�gi�v9Q"`Bf"�I�d����zn�>�S���>9���"DJq�ݳ�pppŧ���;�D���1@�q4���w,��Z|Ļo�c���s��n�������C# ���!_�	�Uff�3X�	M}P�h�����,b+��N��� DZ��B.5;0l8Tj4z4�4 8�H��D @��0�BF21���da��!f&�xF2k�F, "C[U��# :A%#ty�Ð���+�!�8P)�Q��U���:G��IBpޚ�H �<���o����H@�W�S��Q������C���B �C�^��炀h !��"���������E|��_ؼs�J4�RBf�J#A{�C���؆��@x��/ڍQ*��R>\]��f�������  �	=�
r	��D�$y܍Z7�Z���Z�Vجg�\��$�f꛻���l�=J(��}�}��%HъԊtfW�s.�ٖw�?U�􉦓�9e�˿��l��}`��<��U����UK���#�;��� �� ���A#��1�s�~OϿ6H�����"U(`�߷�1֘��)<���;��պ$�\�u�I�ڦX�/�?}_c�bZb���0��#10�q5S�i��FA߽�|F3��-��)T����m�����qZ���dƜ� ɏ�7w���;���/��Iأ�D\G ��C�8t���>���^���RT��$��nt���9��<��� ��߯�����o5��  n��\�E1�����͉��t󥊞p��N�FL��������DW,؞��#��gj�
�ɲ�Lv{6Q�s�6��\;�k<��8㇥�e�cGk��g���������bԅc�fF��,z��jzvrIn�G^R'�
��q�9��������%Y��4��;���	�$�;��7�{F�ˉ9^�l�u%H�@RE|�p�ܿ���o�c�C�8a�+*�FK�f�.�t\Zy82��a��H�N ��e��>T��܃��ۣt8_"��t\Zy�\����l�ZL0� a&�P�.�;��2�>T�oʶt@b	��5"���à�f�]k��j���J�f�x����پ�	�5t[�@^�OrY�  c�B�8K)R�S*T�� /=���&۝1�m�v��N2e*��I%Ο�փ��{~hw�"��sv6�-�3��p�}`���2탸��f�5���c%Ώ�v�l9W>��9��5�(�����^�)�r�svp3Gn.ٺ�]���y���H�՜2�~*��+�;���]!�È���뗳��wI��Z\�d�R�	�H� cև;���8".  ����8 �}���r���r�q���q��������:r�}��>Մ֣�ċ�$��ǈ};8�� c������@��<�~�;g�Ev�����s���ۓb.��iɂ�ݍ��H�za���1C�|0�6ݽg��[����m9�cq�-�=��kج��P��v Dx�K�(R�HD��E�֘oZ`@ �uQ���;7�P�("MM*I�@�ht㘾���H���h������u���se0�a2B�G���nޏ��	徰P~UQ�v&��>�>�{*����V�6�\Q��)����Z<8��J"�)��E)��j�� oϯ��9�e�U4�i%1J�;z�.Cu`�ʹ��<sʓ�7�9$p�l9P�o�g��ը�1C�v�T��E�~����/{�����M6��ȕT�g�� ����C���p�ߞ�G;I6�  �z�R5Ӄ/�����ь�ڷE;WPN�=�һ��u��Gq �{0/��Sn���V�Cs؈�����6]�`Sv]9��m��۷U�'-��A�5v�%A�YiNL���ER���9N�,��-���;qZ͌�-+q��(X������w�����#��-���6�D��S^T8�gyy�ӽ�c�';\�[��v�(ʊUID�cs�ioZ8���B�f# ��Q�-���� ����ƻ����l7*d`�$u��縸6�{ӛ�}`�Z���8�N��ƅ�@]��.��p�Ѥ��SD�/���r\~<�����b(DK,����x{lvf���+9�j���:�Kߛ�|�bɤ*��oZ��{s���Y��\�2�F(crN����@���p���	@ >N����f{'��׭4ۜf*Ti޴-���3��O�^t��3��c%΋�`f\�>Zy���,�`��P�2�����N���B��O��������\�S�d��nNڲ�n��E ��/b&�TT�3A$bRF�rY��7���������!�iȡ�g�9�� su�o���>��'ar'$L����]w��@̒D@� �<���twW��(�IP���H��o�.p��s��qTT����:=��yn؈�Ս6�`��[���h@�q�s`q
`����3<{d�viv.��lV\��߾���[u���ܝ!��9%��UID��\��ːg�O37'�b�f dQ��F��O3=�����v��H1$"RF����3(��g�* �9 �1V;H2� �
LQ%�B��ǻ�A�J�>8�7<�l�Z�o�U���><��4ʰ��m"8털q���c���s�x;��g� ��85@Y���
�E��塽�������(�IT�Ai�[�΃�*yn�ϲ�oi9IR4daG#��ux�ݳ�g�3=�nWKe79�B����HˬSo�W�=�$nC��e��˞�ʼyo��{������ΑI6�n�t��d&C� ��.1��Bz�^��C�ҡ�B!B@��C��eHHA��WU� H��b	�$'��N$��f"E���!:�E'lB�E������\�	$b�4(C&d�D&m/i�㸐��v����тA! ,X� r��0�b�`D �#E�b�$`I �'Af�4��aǨ�$	$$�S����q�7��cv�dڪ  m� H�Iڵ�z��  ��              ׮�r����k?�>����
��dv�>�x�ޤ�R��lc����pF�GkGCl��q��+ԯ4��^��Wn4܅�7�h��ϛa"9���v�*��U��֕qv��:�ʐ=� 1E$̀�*�a梪�U�t��R��%U�B��K���F�lRgn^�R�.6CL�-u]�fU8l���u&�WWl���s��t��<N�� ��!e���S�s��Ű����j�oC�鼗	�@���q�#��̇�{/l�i��1�p�BR��8� y�&��LE�Eq��n.�[��L��Rtk��ݑ˷���	݇)�U
�]�^5�']�`e9�Tx0&��7�N�*��WL�k�!Ul��Y��j�b�&�JۥJ�:v�S��a0�b)�{��5t�����R䰅u�\����\[��\�I��!�K���l��U�����47gR�e�����8��<]���7`.gb�.i��Z�"kls�O ��B�WV�6
�j�I�ͭ'6��ۖЪ��:�ݶ m��	WZ�݀^��,Umƫb凱�ڂݺ"����^f����5 9�Z��J�ZU����0� t�a�-i9�^���DM\�n1�f��F�g��.���"�Ft /T��*�Wj�Kn�i��n����P��յ������<3�q�ѷ�On�q��MlbkT[�kd^N{lR��_Rn�桶��eYW����wc���}��8��ύ��u�t ��@ѷ���0C�~^��~����)��(=��.�?x�����}����8�H�`  &�z�r�Ĳ�{b���X�\��f�Q������37\6�ґ��Z�[N�)*d��4�v�F�;���u��Zw�6]�l�n�j�.�a"s�OWg���r�-l����7E�*D��ˈ�o*��պ8�����<�Hq�G[�.cDѺm��e�6��:T�"�4�9!���K{sړm©�yێ�6�s��"�7�4m��](���I)�$�Q�����nY���ȼڎsp�3TR�)!s����E�g-��g�A���
84��*��F3{���xD�43'��A [>d�4��Jh�x����wb�G���i��r4�`�i�[��zyo��[���܂\��C�v�\hP;��^59�;��Z���_lRjx���Zy�r6��-���X��Nr%%H�f��P* " A��o����  ���{S%)%5D��#g���M���_X>�g�01$�へƎ���,�9��z �-����vR���"RF�n�����E��gN%��B]�)��F۷�h}[fٺ;�yq@40�=c9��s�6���$�'_O7}��n�[��C ��xų��Ji%4dʮFg�@�Fc��y:c0n/bNy��R��D��e�~���:����tD"A�Nn�(w�s	�&R�)TJ���聰 z�0޵d\�����45�(��)@�̴:!�g.��x�nY�,vw ��AX�r�v=��lN�Qn��a�ڟ统��ne�9	}�o�Iw���<ypB\�����D�n8�/���A�T�3�Tv�l��.R�
��I+�8�J#.�_>f{ �������!'"�x����߾��w��<^��E�J �"Z���T� b�A�R	A'�T �Ù��?�����͉�(����5������f{ ��tM��\]2�}¥vj�����+�jJ/g&p�#��#IiUU����kH�u�q�Sn�Cm�.�x�W���������d����J(#������BI�����L��`nd i�Kq�܈���/5��|0;~i���ꖥ4�ܸ�2怼֘�zP�i�s<�'�� ��u��%��\F$��  ��p�3)�s]\+rq�⣷g�������&y�ș۬�.�`�]�iw��Dj݃e�%̶�0�m�*T��7;\mF���� n��W�Z�7�o\�m�gu�2�]*��\�sŁ+7c<�.W��B��+�y�(�-�S�(�9Hl\ݞ����7b� �"�{�w/{�}�>�DͶE�ڰ�^���E���|����b����	��Ţ������o��~(�w�"nfo���椷�%���UBIm
8������8�3e�ѻ�&d�0*ϓ�Kq-��r�3�������������D��[��Z&&k��`fN�2ř�T�=,�9AbH�(�c��_�$��89�n�t��Ϣ3>i�
-}:�D9	���ݐ2 �'O=Ƕ9�ݮƹ�r��v�f(��ށ�NY@ww�J�36X~i�w>�A\�2\$�u�� hp�#��h{�M�D�Ƃ� 2n�>�8�ˇ3.hߚ`]�L�4�.�X��՘7���-P���`{,=�ʼ�STf�D�%�P��q%y�2"̖oZ`_gF~��y�]���ok��9�`Z,��ɻE�H%�GY�F�R�Ȝ�����M�~��:0;z��ك���_>��O@��O�s���7昀��XF���q�*�˝�i�?%\Iu*f��`w�4������i�pӖPD^}I�^d�;z���Q�~��T=Br(����@�o`\wa��֟��ģL7�b���qNָ������*E����Ҏ.��f��d����s�7�4���CןR����,8�GI5g��E�z:I7��'���$�Y�	�\p �1��#��R�
͖o�F���S�Kq-��r�3e��Ƙ��~J����Q��F�9���ٛ���3I�&��7~i��3a�w�ߥ���]�~�㡷b6L��p\z��Lu�M�x�:.���'F���Pp��,I#�|bZ��{l�����2�ZP�z��1-1�9e��0=�4_�`]φ�<BrB�Pt�����V������>֘����\�'2�̹�2����C�`{,Ƭ����Ci�����i��.vX�i�A�#��\I>sD��=>m̦�� �f[  I7l��,��.���(&z�h�*�N�
��"盞	L��;(�8s����념kK�Ҷ�cu������%�x�O�7� ������1��y�����Fj�5C��gm�;�sI��m���7f���Lss�Dm�gt�UwUK��� �1!�7G�7����˙����\.Fm�o�Α����Q���\�$�ص��Ɠ��������w������/'��y��ږ�)�s*�b3},�i�۟�4���h+
N \&��'o����L$���`la��cjT�K�T����Ƙoe��qF_�0=���D�4Ȉ�l��Y|��R�͘p��T���O�p~ತ��F����jbb����{ѝ�d�i�ܱە�!���t�*Œ���Do��/���>>����˜�$�Gs4�����|�������?�Z
�!�B*�Q?_{����HI�`q~�sy�J��]2&�s�HKTl�`nnң��.NC�߼�o�BMD�6P č3�H��A	9v��0�$���`w=sʖ�)�s!@^y��s���T��`_��R�dQ�	�)"@�%1��"��{��#zggmѮR=�N��]�)N[v�I���NkC�D�;D��I��zL��J���P����Ƙ�i�}֟�Q�Xl�KR1�L�㽀�y�A8�j3;ϻ�Ou�)&�m6^�X�P��4%@�p.�>Ny�T2g�4MX�XH.� �p^�� F Bm����
ؤ�(��ĩ)�	�A�[�ˬ�9)�,	 %A��j'"/:���C��D4 ���yF "�  g���>)�� �����*��!�!�/��1���<S�Bt~��w�4`nO��r �@�Kq
T��\�2��n|0/������HjD�\�KT^��ۜﶕy�����ȕ~��
B�%$��i�p�L����ݗlr\Wh"��o�ttN�q8��0����4����ʠ�~���.3�fT�j�1%�֘�[J���L���	���Ԍ9"}�>�>$���nh���	e~0�}�BO���4�A7�&y@e��np`^�LG�*y�Z����ԗ��nH;R5��qZ���0/����Dfq��[p�D���a�ڹv�,70�4m�$�4��R���n����@f�L�4����?D^O��`����q
T�F��i�۝��t�.KY�G ��m�>'�/������cLߚ`vِ7.%�m��y:0/1���Ra���&rC>NeK��H�D�}�0=�$��Ҡ2���>�8�����B\�H"D��
"�(E*� �#
�^I�'ۛ���c�36  t��䈂u��6��sJ�(�Rċ]�'���2;�ڑ�Y��c�����#N
�h�c]n�p
 �.��b-Jm�v��$���͇�[�I���a8��m-v�d�s�F�M�U��Ӫ�6�Ҭ��ۘ9ݔ�s���5��u�d�t��涏�����~�L���8!̻/4��3
S	l�.��cc��h˹�x<�]#��պ� 4���O$9�`w�|`_q�n~���kL�6��ԓ��lt�s�N�ye�a'}�/Q9^��/�ܐt�vp`^bi�ĹĢ/'�/�0-{!��"e���d���nҠ.3a�Ѹ�L�����\9��R�P�`_gnta��m*AQj�"=�M@]�sú�Qɺ]�ǫ>t�M�d�F-L���T�3��,�hGI;_�$����H�9dnC���9�D�[c�������~��\��7��c>�؂�~C�!�'3.�-�I@f�L��0/���=0��;{��$a�&�^�I�.M=1,^,�=�O$s�4�arN& ���@eΌ����Ƙ�؆�w~���~���a�:#On��<��<g�ۍH	�.�iFf@\2"
H��'���A��L�������$���'���A��L*/��ܟ��`o�`��ɗ.eD��3g��83�[\�R�$UOES�����$�}�N���ɹvI�9�l�2���90��Ƙ�сسT`��S2�%y:0/1�nt`_m�@	flkbp��9R��6$��(��\R�G[<��ɨ����;6��\)nbJsZ`v�����ҏ�3g��fәnSmʘ٦�@͟
�zP��w�0;�� �L��Z�$�w1�.t`{�w):����ƙ��9��Pۙey>x��:&%+�\�X��YR�P�0��L��%�f���cL
�zP�ц������v�ؐA��.���R;>�����q���b�`��e��S��	��O��tt�/���I9����?*�u�����ȜiKU؃s_��>x����D�tc�d�m�%��͟D0/1���*�oJ� ��Dz\ʑ�)�c��o��P���Q��0;�mDn@�4�c��]�}��OĜ��;��ɲO�pZ��B@�E�E<@�o���m)�cf�wwwwt ��Iw�Z:]�l�kWZ�L��v&xIw
JQkqa�n�ISa�&&Q���ڑ�n�KtGn�pV��];����p�f�]��n�V8��+��n{%���v�mѶ�;Gݵ�3�i�+pS�<x6�KW���y���R�2CE���N2Ɠ�0��:zd�/?����{��k��x�KjMI,������SnLf��oR��T6�nm����9�J%��nZ�7>����N[�G�`��-;��cfF��(���$��d�y�����f��%6K�66P�4���#�o�y:030�S�ܶ��T"u��D��L�ۭ(���S��D�^�q��|��ۃ���~=$��L$�0=��T�/���˖�1*X�Ok#���o֟O�����lv��R{k�󻗞��hl�MD�`��`onҠ>ŭg*���w_��9g����@|@p���MI������i^��}Q�� �Q��o�<zI�f��#|�Τn���������p&��;� ��x�/g���oS>�LF���9��P��@w'����ݥ@_��D忺:I���^�DKH$"E8���<w=Ǜ�s� �v���fK���_|�ˢ-�uo��4��cL6/2�Wb�#g�un�I)�#���'=���$r�t�R;��n��%r]q��|�F�pt�wf�o)�~ Ę	�mI��\vW���%����[(>J3_�UL��;�~J/3��~#�ܩp�"�1%��0>��Ң�/3Ԩ���$s��l4��#��TEK�^��t�;��V��[V�iB��8;�;��q8�%��w�0;w��q��Y�0;��N(��KPL��6�|��\�7����y�o�6>�7Q,s#r��-�6|0/,Ԁ�Y}$���'�N�&ˀ���l��8����R�/5�n�J��R�����!=@03��ɲ}~���$���pt���'�#��-߇ě���[$����I��'i�Is��;9�y��X�ݞ#hiG]����w���XGu1"%�����@^N��k�$�@^y4��/-ю%���-P���qq#��	9}$�-��� ^j��+�0�5
[����4���L�r#�ݥ@f�9i����q�J1�K� s�_}I����P�����I�~�0�uD��KPL�ٻJ����k�y�"N��Y���t�I��ۦ� ���"�0���E����"@ � �"D�C���/^�� Ha&��Jd���c9$�<@��A�|z�(��,$R�$ �aQ}��l<;�.�`�D�F$I�Հ�DhE�7���FB� He�a#J�2�zހ�ł5"2#*B*��f �#�G '��)
L D �(S
B �M��-�|�� m�8E$��b�8qoS�C� [@              m��j���2�Cl�����f�H�e��^���M��v4X�.
ڸ�{e�˫k`m�%7tZ�Y�V�����F7��M�GF�\��퍀�Ά�l��.Ӳ��2�AŜ�[�+2Fg��6l<C�ml/%ҫ�&vƒyI6�Lm����m��Q�B^yյ�Zv�'+Zn��TϯD��R�vӨ�1�N�v���E:�ᣄ:�b�s���{=]/I+��8�nܑV������]���mb������XZ�@�r-4��҈mִnI��	g
�;7"�jܞ���m�mi���6�Y:� ��,ƫP�4r=��=,K��&�X��6����k���l�G!UEfz;K���[#i�iZWc���a��[%�yƕ.��Ƙ8�6ɓ��dݑv�^]�8�%[k%{X*M��p1�,��{-��K��G.�:˭�b�4ʈ�W)h�7WX]me{t�ڳ���ë�m���s+$fћc2���djU���D��u�^�V��AUJ�����c���h��-�v�[��k(Ԗ*.N�-р"^���JKW ҷm��� 6ٶ�� Q�VT���&ɢu��rQղ��U;�"���mpnÝ[T��"��H
F�n]֣uH-�܊���*�ʫ!2c��1vd�C�>��dXPˡu=�������b8�	�족\��Ԇk1«�NsS�(q�u��N��$U����+��,�&��'<��?�$�T)"�� ��O�� ~�Q��Tܠ?c�T8��@�B���Do��%@����ݴ̛if�wwt =f�B�����7;j�m;l�&^T�rKf,i�,i�����6�(��\�B���,粗;%�b}�m�.6r1��lvts�n�ݼ��WI���ɣ0��s�2�Z�lY9�Υ�\��k���cX�L��dVŊQ�j�Η�h��z�!&	+��>��������-���'f9籸��С�.|�rے�GhD)i�O����%�T�
6��=�������!��'[|=�ץ�R�K&(��*�Z`z�)P��sARJqH䁇�D����w��^O�n�`_f�\��8M�D�A����Tv#6|1�4�"�Ԙ��1ĲSm��T��a��L�4���R��1�"93���4fG���iSF4dmi��C�3�#�|�c�b�G~v߽Ђ$��I��po��%�x�M�i��n)a����7}�@�^x	�%$
�|V*����η��&}��N@�����c&&uL7�Z�ePllk�@^N��i��֘^"[���(r7jF���]�!'/��&���=$��k�*%��-��7Z`Oo)POs&��r�3�X�[9�(�Ɯ���	�����mӼ���	�⚹n�o�`v��@^O���7Z`}���r��p��K]7_�y:0/1�oZ`T-Y�K%6ڙl�/'F~y��/�4O���)z�>��d�]�(��F̹M̒���(�i��Ƙ�zP�����.�*b!ʠ/5���ӠfφlFn���du��c�np�Sqk��N$q&wu���S='E�7<=�+�ʑ�S�.[$�Ǥ��L'���:���!'�M�\�
H�=!y>��3u��`v�����@}��ٚH*�U��$＂$�4��
���~���j�h%�m���=m�8I�֞o+������(�����^������6��Zm�1����@^N�	��Tz=7��	���>͞�?6CIi���Z\���Ыۏ]9.c�ᶺ/��wq�}�����Zߜ��`^cL��0;v��D����l�A%F�%SG����� ؀ �'�$�������3�G�h���R8�IITo�D����s�rg6~�i���R�MHB�"��'-�=$�za'-��888�|��%Șq��ne��l�`f�Lߚ`v���4AWD ��I �e��ws�a�M��  �wHV�6j�#ѧ�O*���c&U�wV�e��8ͨ��6��7g�Nӹ�w���N��t�Cgn�`�G���#�ջ\�ۇ�����iΩL�$.�$��Ď�r�H=�b�)wTs��v獱�)l��ە��盈6�v�.̏5��s��3�������{�w�o�9�,�ɮN�glR鱋O4{Jvi箈�@���p�l���0;x��o��_$��ƒ�?�|����	r9 n�r��~� Dɼ��	8�J$�b	�� DU�{Р�(��i8:I�z~=�F��%��$���z��6S-��M�O������־�ϚdD^c��;��h7	�jy-�I@f�L�9ĕ�Ҡ/1��/'����'2�B� D��ѻ �x�]�.��z�$Ӭ �OI�s`Jg�|����b���\K��q.�o�F}����-�C�ʣb3u�W�s�� "��Q'Gui�&��J�
���-R�*[���P�ၹ�J��0;v�P�gf"%KR�F�%���y�0;v�VD#&|03'��Kr�R�@{7Ԩ��Y���>������MDC�J�	��A�Ϟ�P�۶���SB-v7z��,�$��B����ڀ��yqT�`w�P�(�HPI!T��s8�J� �/kJ<�����y��<�@ U�|���T�1%�O�o6���s�!W/��G�?������Q*7.T���R�Q�������a�㟷��@w�d��Ĺb�(��������@w�7k�C��~7Z`_�(���Ie��������]�ѧ�j�t�L&�c=s��8Pۙey>�����R��~(������pȉ(�i�ĒQ�+�BN[<zI�ǌ�8��z���!�m��7�0ؼ�Ҁ͟�i�}�d��[���	j���ݯ
�͟��;��6O�`�$Y!څ%�b4"� g50��\��)R$�[(���%����4����A6��"(\D�e�	�
(��)v��\u�n��n���1"�2	�2��I7v	��$����8�%�G�'��hߢL�ܹS�h ��L
��TFzx�� @���tv��T�J$�G���T��x���0/efMȔ�JARC���.��$�h"Mޠ��s�E�}�@�O�T�j\!��P\㠂$�@ 7�'������/҉��������?}˛�iL����  �޻�}�����U���TK��B��۶1+�@l2)Z͕����G�.f��A��y�M�h�b�n%�;=�h5ڢ�{i�i�Aw)tm�zyG/<{c����%\�u[r%��')��ʵnm�;����5'nQ���ɘJ������m��P� �i�o]l��\�2�,�g>s'ݜsiN��V����K����u���^r��^�kL��*#6?.q$�7Z``�?k1&�<2F��wZ7w��I:���ߚ~�\K�ayf�7,%9mL�T��lf�&��[�R�/3�TrC��cjT8C��3u�ٛJ���R�����F���Ӊ�˕1�P�i�ۼ�@df�^cL�,��B]���p�,�b!�6����F;ChӬy�J�gl�Woǻ���~~+Vr��ߍ�ݞ=$�uLH�`��[�!=W�]&ܳw���9$�����x�)ؤ�@���B
��EB����5� �>� �=�L��2O�kI�B�K�4ۊ� �ﾥB�i��ĔE�?��N��E���!���pt�o���ݬSó.^�'�@�7�s)���a����y���.qql�֘~i�Y�Dc�.Z�*e0�>��a��VO韾� �m��:�[S��vݹ���;Ke�x^�����Py�㣈�d���È��I�v	�p$m�;�N[<zIվP��8+�aIa��$�j�۵���@�tҿώ�A$�nۖ����i���@@��aU�ڝ'I�H�(3)Tj�ǣN0�HJ�ɷ�C�t�{ �f�t1ނ��f�gI�#�i8$`<*�U�<@8��s���O��R��1�������q�c��������̇��ߍ,����$LA �$R
	
�̔�e͹.IR�N�00�!B!SS0�`�_����%�¸�̇J!�:�?�@�(qj���i��?� ��| ���w�����A	=���N8�rL���yiN���P�}�i�w�L�A�PJ��BRUH��N��	>�7���7�9�"�ϧư!�p��fu�wdT4t���v��N�g�n�0Ij.��nh��֘���oOs�"��CԨ��	N2�s���N�{���7vx���|��݂w���0�h���5@f��@d^�^cL�i�P�e(��9C�}��|�&��	���'�;P{P�;|+�3��NH]�{ÙL�J���3u��4���ҀȽ��+��*bu0��%8E�n�lg�t��h��M<-t��b�����_Y�a:b�3MZ�|��oE@d_���ƘNk�SQ8�e�)�|���ǿs� "���	7vI�X!'<Š�� �7�&�����C�9�����	9��P�kT�R�7�n(>\J7ޤ��֘�~(q�\K����z5�a�H�/�Z�3���s���V�c=&�D���z�kR���*fRI  :�.��.�6�m����;n͒�B�Y̃"l�������vqe�bLv��ܬ;'k�vM��� ��c5����u���&B�Rad�nx�y;"y��{sqev��v3�<t�뱈	�[]��^ �RY-�Gn�5���pMw3[;:nȊ��d]��;���je�{w$\)�99��Rۅ��Eܛ��&~\\\�U*0�Hm�t}��P���Ƙ���wCq-��2�@d^���r��7�*L��� #�d����nn���n^@�����0ȼ���63�ɏ���~((�h4�c���/~�D$�OI5g�D��!&����N8Cn�c�/1���(\����z(�i�~Ƙ�=w��%	,4�@����!�t(mi�ق�������i�21���'U򄜸���}Ī�7k��_z�J�,S($���m3φ�0 )�2�2I�zi�&����[����i�8�}���oQ�%�(���0)m�*�}��ĨiC���z��nQ&�D興���ٽ%���Pܵ0�@d_���}�T��l^g�Tf�j#�	�@G$�)s�rFDğ4�
m��;#b+�L�q�2aƈQ�ĝ�����J_f{���"u_)ԏ�ѯ��JeDD9T��P�m*c2�j{� ��u�N!�
���M��GN̹{!���z�Ђ$���~���e�L�(�������CԮ��}�0�s�/2�(���2�7�n(݂r�'�[<zI�|�'���*�z�n��hKIo�'c������1�B�G��{�����|���|rՁ�i�ۼ��2/�`^cO���e�(m�P��V��2�6xI�r�rI�h/d���H�@܇��W��?���``Vc�Ey!�.T�rD�����0/1�]�(1s�~�$�s��Ӌ{� %��}v|T�JJ"���z��8��Zt��0.��8~��l	FHe2�	#H�\i��<�u���S<�����!a2�e�)��(�����Ǥ��r�>1�x�v�~�%��zR�nT6�S(؍������0*�i���$}�<$H����(����v�&��;����_(I�%(6�#M'j��kL
�xP���Ff�`]ϡj�!Ķ��@w1��.3a�y�"Om��?"`D3��R�E*�u��  �7nٵ��v7ӣx�4J�k�0�+uV�J�8,�X�c�LkN˕�Ԍl��]M\r�tL� �-���c�t�m�hب�a�m��3�g�����uŷVؕٛ���`67贓f�K��DYԔ���ˍ�nMؤ��B�@�]j�Uh2��.8�]��a���V:A���3o^�̓k��]��gg�����n��m�hx���ĸ�i�}󑇣���f�=�mʗ0Bp9�o����0;v�zI�uO$~���m�N1M��q�I�����D�K��N6�>���h�R�"&�*�	�Ow�<$��J53y�0*�|`^��d���8�.3a��X���0;v��3T���4ɭ�+;(����j���tƎN�h�0�]����,c=�	�Je�!��p㽈7�i�y��w'�I8��$�d�6�#m9���'ؽ_�%�����zoz�P��i��ϲP�Gq-��To��#}��Ȍ�4����B��bn�8�"Y[Is�q$�_��%��T��0*��P�D{B�,�1@{wԨ��G`@�{��M��x���J$��s���x6x�q%��ѱ����ӝF�z���Q�g�dm��8�l|A&��	=̔������I�`q��cN�!7	*>�]��^\\�"��035����"7<5��p8s$9s,��`fcL��~G��fD�?E+؈���Q�K�`_�~(ۯBe�!��n(݂$��+��[{��M[�	9rR�s����U!�Nf��>�"=  �t�'�ߔԎ��	3�\�~��P�܇W^ƞl�m�P�v5d����s�e�Oa��f+�w3Ԩ��`fc^\I.%P���D��x�'j8N�uo���i�.����ҾIqD���ܗ"m��D�ނm�!�9�p�����C��)�ˉ��$�Po9���"Nf&xI�͔O����0�! ������f�l��w�r��r���I6���MWT$�`�H���!�hp�\Jc�l����c�����OF�JR�&ӧ��]��<�-���������֘~kR�*3�����D��p4ۊ�A���f�����P_)�8 HݳJm�F�nqH:I���xQ��`n�L�~r���Ħ�D���IF���������֥��@��Љ9!�	M*U*�3H𓓟C��0�fz���?�#�=��A$�nۖȨ�ȑ���1"H�1![[!H�РH��B�$=W���u �� 	&��I�U+ OH�$��"yM� CC��ĉ�� �(�+� D�t���")�(~N�
�k
����|XR�  ���_n���pA�$<�;�vo��    -�H��ă��8$8 �               N�mѮԪ�N�G�#�%���vNOn/[-�Wp�G��]D��>n�T2�ۻ	Xכ�#i�J2Bqvz���v�Ÿ.�e����v�����U*ܛ���*U���掉�YY8Cj����Z5#cd��q)�蛒��֍�h���9˱�5XԙzZ�ۮD�ɳ�U��Ԏ]���1������ݢ�����gvȫ��6�)B���䍹V�!��r��4��1q-�Wu�S�'F[d�i��q�-+.,ڻ9���	��u��\�\Q�`];�pkp�`�2 ��epJ^�uLm�ڴ`wi;�jΌ��P�u�u�{�u�y� C���M��\���ٲ�O�j��P`6ӯL��n�ѱ.�A͉��Ǎւ����m���֣n#/\zwW��Om�p�[1��\�yS���<�����!��[�YƻL��ղXr�\5��`�=q��.�p�{
c�YmK�a�ٕjU���-���N��2{l�[�m�*΋h�&�ćQ��gX��`%�)V�fl�N���T���+Oh�V�mT�U^U�X��
RZ�YU����S�ʂ7s(g]�zb���ι�����Ch�ೲ㬎%ئ�uڜ�[2K�(��*���iT]���l��.��A��6�uEs�����6k,*z�L�/e���b��un�Y�%j��R��u�� FX��/6�[cq��X�-��e�݌݆ᛓrDE�<�P{R�$W�O��J���G�P$ �s�`mU]$�UPB�5��  ������r^�|]lK�<i�6�&�K8uz��QNs�mb:����n�F!ݐ�݃��ރ�z��u�ۉ P���!nG�.��S����iwt[x2�n�WY8]!�J&U�vƕ9㴜�������^+�m�{	�jË�K3u�>���x�1���7\y{']�������t��uН<�X\����;�v�ΰN�����x�@w��Iq/�8��z=�0���Q�nq��$���~�%=$�|�'�`�#o���MA
nceP���f���0.�����
��q¤]'�׾P����+\L>\Qv�ؠ=�?J%>C���P�i�w�0;�܊#6�ؼ@�%yC3s�{�g8�v�ᴥ���f-bk�ў���{��M��*q�;�'w�CԳ7GGI:����U�֘��r���r؈j����τ�*��\��A7��y$�b�ď�g�tH���8:Iվn{kL�z�w�@v���2�!���֘x�G{{J�ˑs��pGl�쪔���Ur��t�ޠ�?�.��]c~�s`_�C�4��9r�܅����F��D�.崶��c���Q�d��q�"et��*#6�i�w�0/f���Q�.:I��p���BOsPD���6d��4UAB��S�̜��d���xl����H)B"D �T�����N@�B�:Mt{���\ߥs��"�AJ�D�%��n�D��󃄓m�'��Vn�07gc�%�(��w�R�ݗ$��4߂ı,N����"X�%�QNy-�Ep%��h�a��i�'FܕZ��Ӄ-���YL���O���iq�{��g��%��S��dK��}�Ȗ%�bu��4?'Q2%�by翝N�X�%��p��fl˦��'Q,K���jr%�bX�y�ND�,K������Kı/�}���bX6']�=��]ۗ6C2�É�Kı;����bX�'}��G��?��2&D��~f�"X�%���p��Kı:�=���雙�It�uı,O<���Kı/�}���bX�'~��S�,K�~����ב9��ș�2%���l��%ݙeٗM����%�bX���٩Ȗ%�`��5<�D�,N����bX�%�>�'Q,K����
2xC�.3 ,�a�0�nM�7���6�v.;1����=zC���w�{��7���>���"X�%�N���5:�bX��|�Ϸ��Kı/�}���`ؖ'�y���f�]d����%�bw��59ı,K�~{�N�X�%�|����KİN����"~
�TȖ'����sm.�ٲ\8�D�,K��ߛ��%�bX�Ͼ�ND��!�2'�}�S�,K������bX�'Xv~{&��ۻ�d����%�bX��ϳS�,K���xjr%�bX�y�N���,ɑ3�{��N�X�%�৿r_�n�fl˻%��uı,O>���"X�%��G�~���%�bX��=��'Q,Kľ~}���bX�'��E�����fһ�6m�ww@ ��I�N;,t���k�nUn�Ƭ,���f�u�	c����{@��$�=r�W�鱹��v�K�Ayu�wPmS�#�d�q����!�5���[��mb�m��f�k��3������Y�����ZV���;�G]'\]��&B���i��%�B�2OL�{S{������?u��f�c[r]�>�a�O�smU��#x.�͊1Yu-�(O~����,K���59ı,K�~{�N�X�%�}�}���bX�'~��S�,K����ۗr]3s7t�uı,K���N�X�%�}����Kı;����bX�'���S�?l��,O6�O���Mɦ���uı,K���jr%�bX���ND��a�2'�~p��Kı/�{��N�X�%����>�2f�n\ͻ��N�X�%���p��Kı<����bX�%�>�'Q,Kľ��jr%�b\��t{fL�ne�ɚq;�bX�'�}�S�,K�L��y�w��Kı/~���:�bX�'�}�S�,K��Q�����ۢf��TJ����`qŻS^{=��[�GX]�l�6�&f�\:N�X��}����uı,K��f�"X�%�߾��9İ�����S�,K���>&��ۻ������%�b_>�59�������W��<�bo�59ı,N��"X��%�?7��Kı<��\�!���ٗM��N�ؖ%���p��Kı<����`ؖ%�>�'Q,Kľ��jr%�`؝w<�/Yvfm�f[�q:�bX�'~��S�,K������%�bX�Ͼ�ND�,K�}�Ȗ%�bu��fnK�.ݬ�q:�bX�'��ϧ��%�`�߾�ND�,K�<�Ȝ�bX�'���59ı,N��ލ��e�1���V�㓎^�#�ּ��Ž�d�q*OT��3k�ل7&��l8�D�lK����Ȗ%�bu�59ı,O;���"X�%���s���%�bX�}���sd7-�����ı,N����"�ؖ%��~���Kı>��{8�A�,K��٩ȟ���,O|��K�&k7.f�t�uı,O���Ȗ%�b{��q:�c� xt��zh>��g ؗ?_��Ȗ'�S"y����bX�'�o���sc74�]8�D�,F���~:�uı,K��f�"X�%�מp��K���ϸjr%�bX�&�>.��ۻ���o��%�b_>�59ı,N����"X�%�ןp��Kı>��z�uı,K���I~�e��f�o�.�m�~Y.{\h��4�N�^X?������vY1t/��Kı<����bX�'^{�S�,K����z�uı,K��f�"X�%��s�r���͹L�wQ,K��ϸ�r��H��纜�H$��D�I����?a�dK�}���ܗrݛYt�uı,OϾ�θ�D�)ľ��jr%�bX���NA�,K���Ȗ%�by����wr[�\��N�X�~D2&}�����bX�'~�xjr%�bX�w��S�,K�*~���7�3��q:�bX�'�����wHn[�����%�bX���ND�,K���Ȗ%�b}��q:�bX�%��S�,K��(����_��.i��nvn\��'��\";���z�� E�����]��R��w�%�bX�{��S�,K���9�N�X�%�}��5?'Q2%���=��NA�,K��I��l&��.�N�X�%����q:�bX�%��S�,K���<�bX�'���S�,K�����3v鹻.��uı,K�����İ��"X�%��s&�"X�%��r{x�D�lK�}��d��fl˦��'Q,K����r%�bX�w�ND�/�r'�s���"�ؗ߾�ND�,K����.�ͻL2�É�Kı=����bX�'}��'Q,Kľ��jr%�bX�{�ND�,K��������u��E{h��-�  OF�aa��K�uΤ%."��g$��8#U��t�S���9�����	�����ڪv��o���8�8��/���0V���s�
o���Y��GeY�����Yl;�3��s�/N6�B��]l;P=;U��	l���n���т9u<��p��%�Ɲ��;!�-��:���狐�G��Y�QW36�0����K3B];O"X�%�����^'Q,Kľ��jr%�bX�{�D�/U2'��=�N�X�%���g����!�6l����Kı/�}���bX�^��S�,K��jp�bX�'}���'Q?`S*dK�������wws8�D�,K�����bX�'���S�,~DH�d�����uı,K���jr%�bX���=�3Y��K�q:�bX�'�~p��Kı;�}��:�bX6%��S�,K���xjr%�bX�'�|��K��ni��q:�bX�'�o�^'Q,K��`��~���Kı;����bX�'��p��K�G�����
@F�
���d��=���l�]�>h)��ջs�9�Θ�{��g��u�}����Kı:����bX�'���S�,K������%�bXr�_�)��-Fc�w����<�g�p��?c=�7�<�@��D�9�Ϲ����%�b}��}x�D�,��٩ȟ�P2�D�|�{�^���۴ɒ�N�X�%����59ı,N��}�N�X�%�}��]NA�,K�}�Ȗ%�bu�/ٻ.d�4%Ӊ�K�@,O<߾�N�X�%�}����Kı:��z8�D�,�dO�����Kı>�l����0�vnۻx�D�,K���jr%�bX�{�ND�,K���Ȗ%�bw����uı,O~4��6nn�sK�h
��Wci�n�9:ZnƮ{5s�Dc�w��.���+�v����'Q,K���jr%�bX�w�ND�,K���o��%�b_~�59ı,O{�}��k72�sN'Q,��ϸjr	bX�'}��q:�bX�%��S�,K��xjr
�bX=�It�M��]8�D�,K�7��*dL�b_~�(0$��>|=�i�m���L	 ��y��)�uu�BH, ��K��\`3�N`D�:6Yϡ�)�Y�.��ó
�[ZXP!�b�hD#�B4�B+H�:@�T�d��w^�9�9��jAn��t
-��`���L����L @�/N����z�
�b�N������ =�W�>M/h�E�*x��l���	��B��;������Kı?;��Ȗ%�b|�S�-H�p"�ǁx�[�٩Ȗ%�bu�59ı,O;���"X�X���{x�D�S"dO=��d��s6e�ng���bX���ND�,K���Ȗ%�bw���q:�bX�%�����Kı?J���}ݺ6_c�;c�[�&ǆ[�n'k\=��`Z�z���6�
�h4ې}���x����Ȗ%�bw߼�q:�bX�%�����R#�L�bX���ND�S"dL��?L�dQ-"Z�.�PqA�g���Kı/�}���bX�'^��S�,K��jrbX�'�����v�Y�7n��'Q,Kľ��jr%�bX�{�ND�,K���Ȗ%�bw���q:�bX�'��9�˗t��7ws8�D�,�H��΍ND�,K�>�Ȗ%�bw��/���K���pC�C�w��~�S�,K���7��ff�n]34�uı,O|���"X�%��~����%�bX�߾�ND�,K�}�Ȗ%�btw��?u�@��F�+�us�v�Y�V��r;��)Ik.�i���{��'���{�_o�^'Q,Kľ��jr%�bX�{�ND�,K���Ȗ%�bu�~O�͙ws74�ͼN�X�%�}����K��:����bX�'���S�,K�������%�bX�>}�'Y�ܷ4�s��Kı;����bX�'���S�.�ș���o��%�b_~�59ı,N���z�fn�a�.n�N�X�%��p��Kı<�|��:�bX�%��S�,K�ܽ���x��e~l��)����Kı=�}��:�`ؖ��s�����%�L��>����bX�']�p��Kı?G�:��	�ӽ��I��_�ߨۋ\�M��  ��\����VӪ\b�Sb˰��	�c��[�SG7\;,k6p�݆ܛ
��;9�v�CH��li;N�5A�]�=�Y��q��N����^�+�N�5��vk�����g�µ!c�I����d��ے�]�ە�{��]�^�˳�#�'0G���O�a�o:6M�͸�ۻ!��/<�wg�\i�!Y�5����\2hI�?���%�b_ןf�"X�%��~p��Kı<��"X�%��}�8�D�,K�~��e˺K6Cww3��Kı>����bX�'^{�S�lK��>���uİ<�3�S�,K�����0�5�r�LӉ�Kı;����bX�'�����bX�Ͼ��Q2%�b{�p��Kİ{�<��&��]7$�8�D�,K���q:�bX������Kı=����bX�'���S�,K��$���.ۛ���N�X�%�}����Kı ��8jr%�bX�w�ND�,K���s��Kı:������f6���vO� �V���ӝ<�Xy�J���$�M�ܷI7oI�Kı;����bX�'}��G�,K��>���y;��,K���S�,K���,�ٛ��e˛����bX�y�NC�pr'� ��B��;�����g��%�b~g��ND�,K�z���g�x-2�͓e8s�N�X�%��}����%�bX�g�]ND����wSb}����Kı��<�#����M�S��!����%�X����S�,K���/ND�,K����%�bX�g�f��qA�X���ba�@��yx�D�,K�}�Ȗ%�v���F�Q,K��>���uı,O�ﮧ"X�%�N�/��l��Rfe�Թݍ8�'n�2v���1����韽�����<�Н3N'Q,K��ϸjr%�bX�g���N�X�%��}���u"X�'���S�,K��=���ݥ�wY�q:�bX�'�������$r&D�?3���r%�bX�}�ND�,K��8jr'�2&D�;�=�~�2�fn���%�b~g��tyı,O}�"X���Ȫj!�;��L�����uı,N����8�A�,K��~����n�n�'Q,K���xjr%�bX=w�ND�,K���s��Kı>�~���b^�dKbߚ0�#a����x�G�e���Kı|�=�8�D�,K���Ȗ%�b{�59ı,O�;��n���[�zl������
b�����u=�o6k�dݙ����s]�s��%�bX�gߟ���%�bX�g�]ND�,K�|�Ȗ%�b^��59ı,O���\ܵ��.\��'Q,K��=��r-�H�'���g��%�b^��59�DȞ�{�N�X�%���N}2��%�&�ܼN�d���xh�%�bX��<�ND�,K���s��Kı>�~���bX���ٙ&hM̻fi��%�g�12&y��jr%�bX����N�X��b~g�]ND�,Ѡ��Ah=�����G� �D�N�~g�ND�,K��4pD�� m�a\]8�⃊-�ߦ���%�b}��u9��,O}���"X�%��p��Kı/s���M�O%�[�<��l�)����'�[�C�K�hHB���M�2�\���wı,O����r%�bX���ND�,K��8jr%�bX�y�}/��ʙ���{�C���n[�n�'Q,K���xjs��"X�߼59ı,O<�N'Q,K��>��S�2%�byߗ޲۲��a��7'Q,K��ϸjr%�bX�w�=�N�X��ș�??.�"X��b}��592�D�<�o�/�[�%�	�q:�bX�'�{����%�bX�g�]ND�,K�=�Ȗ%��̉矝��bX�%'�ߤ��,.�ܙ�8�D�,K�>���uı,O����"X�%��~p��Kı<��}8�D�,K�=�xD�~�����܍�  [z��>��7KͲ�6��v�\�a��#�m�Ζ]�2 泲n��p��\�-0`���^���TT6��ɹ痓jt�h����9*硓��Wʺ�Ag)�W9�eQB�!\u[r$Mi�O1<��M]��׊X)� "E`��r[]��bGs��m�{����y+���.�q�����=�{A����n��8⭕�^�	����ȕۈ�wr��D�,K����Ȗ%�bw߼59ı,O;��uı,O�Ȗ%�b{���at&�ݙ���%�by��59�r&D�=��}8�D�,K�??.�"X�%�����Kı<�|��l���v䛸q:�bX�'�o�^'Q,KĿ}�jr%�bX���ND�,K��䚜�bX�'Fxy�Wm��fm�uĳ�#��٩�Kı>����bX�'}��S�,K�<�}x�D�,Kϡ��ѹ���7s��K�,O����"X�%��~���Kı<�|��:�bX�%��S�lK���vA� P�a<p@�/�6
RV�C�����ֹ�r4��I�j^Tg��~7���{��y>�Ȗ%�by����uı,K��f�"X�%ʞ��F�Q,K�Ze/͕*C���ǁx��7׉�"�x����,O���h�%ڙ"}��59ı,N���Ȗ%�b~g��Isr]�.K�x�D�,Kߧ���Kı=����bX�'}��S�,K��9��uı,O����.]�]�nSx�D�,K�~�Ȗ%�bw߼59ı,O;�N'Q,K��﹩Ȗ%�b{���at��˹3N'Q,K��ϸjr%�b؞w�=�N�X�%����jr%�bX���ND�,K�ݿ_wa�g����\�;N�
�ۦ�ڠ�goW/&nT����w$�Ӊ�Kı=��}'Q,K��﹩Ȗ%"X���!�$O;�`�	�|<���)�����8$�H�{�&��%�by�59ı,N����"X�%�������bX�'�C߲�s&�]����%�bX���ND�,K���Ȗ?����
��� �*�؊��� ��<���tq:�bX�%�����Kı;��r��fn��.\�8�D�,K�>�Ȗ%�b{�����Kĳ�???3S��%��r'�}ѩȖ%�b{��f~Lɛ2]��Ӊ�Kı?>��'Q,Kľ�>�ND�,K���MND�,K���Ȗ%�bw���nf�.��>y�:u��/k9�n����z������5�f�6B˹�&f�'Q,KĿ}�jr%�bX���ND�,K���'"X�%��~s���%�bX�}�Ϧ\��7-����uı/U>��N��DGblK�}�Ȗ%�b{���N�X�%�}��59ı,O|�=�%Й���8�D�,K�>�Ȗ%�byߜ�q:�bX�%��S�,K���xjr%�bX�������m��.���%�`bzy�>�N�X�%�|����Kı=����bX��Q`jT9�O��Ԛ��bX�'�|y�7p�m�7Iwg��%�b_?^�"^Tș�=�Ȗ%�b=��pt�#����Ǹ������3���Z;�axf�׋v�W3���6:u僖�C��K������p02��ޟ.}��c$���$����(�A��'��@.��@�,�i�vM��$2H�|dJ�31�@�,��Q��ٍ2O�AN2�Q��p��}k��h��m0.��@nbzLL6�Ɇۙ�7u�]�Ϣ31��n�6�/ki�m��l�&1 �v3��x�|߽b�TOX�����%,���>��P0Ч<oX�ځÔ�D�@�B0�ؤC�R����4�'��D�4�]�j�u ���z����%�(^���$�,��O׾�>}     ���lHoS�@ �               Nk5�����r�{5��.%���;0DI�I���:��;�L��͵�=g�7r ��U-���4�ړG96Ɔ�'m���;���\�6��UN
�V�\��{]��J*�UÞ�&4��k]�m�\S;,ʇ�Ju�����J���_g�R��yquR�v��Wc�N�^j�Ԏ^
�p�m�cݒv�ױ���vWg�����qH����P��nM��;(m�Or.��8�L�Ib'j�tW�ts�v�}d���+��UT���n����q�6��1�p3�5�ft8�U��V�[�����
�EC�V��1U���ey*�х�wPS,�6l�m"J�TԹ`��p��52@�/�7@� iUs���f�������v�s�k�۳��"4�U��Բn�yoK��è����2������b��kp�3�8�ݚ����6�Q��@3�[�ݬu�[<:��ۄI8��<K�7Bs�撊���ڨ�,��A���� Ά��ʷUA�J�@]6ݩZ����Ug�2���*��e�6X�um\�*덁8�Vɼ�UUW*�삮�JKZʑm-�M�!��M�&�8�l��=Z�r����AX��7+�=�mI����C�j=DL��6��L�S2j�t��������rr/@	%Y�'��V� �w.z��=�Q�.�$jy-�M��s�g��-UAvii��U��ÚX :�7l]:���yݚ��M�n�ٓ��ȷw�~�{��D��jh��"?)�">�=�DSֈ,�Aw�6�H/f����y�~����١b�  ^�7�E����,.x'���7W`ݢ��o�������u�n+���c��ܒh�a�q���*��#�ky�o�Em��j&l�����A�^N��Wn{:6�e�c��<��=��8k�k�Pㇰm*���F�v����j5�7�Vća�m,�4��'�"�9o/Z黛�e�	�L������qʩp�Q�(.��9�������k�:2׀������� ~̖f4��[Y�Zqd]w_� ��`fcL%ݠ��Fİ��R�$&iO����ƙ�%�.D}��3�ַiĎ��L49�w6���03-�A'mp��.���Ia��c�O��a%���@=�;�P������@�n�c�8뭽�,g��۞��ouOgWl&��ΎQ,�ɉ|qP��P�K3`WgFř��r@�ˉ��P�5�_�����" v���$��I���Ϣ  ���Ŧ�F��7����9	?|�%��Ǥ�t�	?[{a�£25�;s�������Ƙ�W8&Zs�Y�31�@�,�i�]�K�_9��O���p�����p��C���ۛ���a�C9��c���壧\��o�ps��_�q#�p��(�~�A�p����k�?p(����/-������̼�×)�%2�3�^φ]�(��b^�s�d���7g��O�fHdľ���c���p����za'U9AN2�Q��l�ݖ�$�Ř��2���ߊ��s�����ڭŲKdX�'`���@)7cQ��U�I�P@Bl&FМ�6���:0/���ޔ����fP�TC��Թ(��+�IDX֔���=���.b�-9��ԶP�zPn����s��:���N!���Py(�o�}�$���~r��y.��8 U���� v/� �o�����m8R�&Y0��f�˝���W�J��f���2�6��ʉ&ͮ$�[%�2��di9�;yV�H���@=Q<��nt}�;yT�7g���:0/&=������"@w۴��Ĕ@o�,�хE��`z2��D�6� ��t���$��7'}�J��h�&FЙ0ܹ��t`;���R�ݖe�9����!����˝���7e���zP�%�_�����~ �7$H6dl&�m�  Ӛ�����ץ�.�m؊8�.ً���iq�I�z�O,�����>����r��6x�Qg����� �����ȝv��f�c���w(O�q\�5TN՜ᴙ �(�Û@8v�kAd#8̍YǞ
9�p��帹D��B�u�^pѰ�lR�7J�S�9w�[v܄̲˸B܂������u`^���n���\Ms��S�'����ҹ@�,
��<�N�:0�qF)���a8��s-P�������`V�R�:��⍧6����4nt`U�
��T{����)�iˇ
be�(�����R�ݖ�J;�v(ُy�BLK�K(��T�#=�;���}��Z�x�D�� �cN<���S�gv�m\i,��nڱ�gÖ#a�ƕ̍�@ݖ\������U؃wGH��2a�q3@w'G�uq$��s�)�с��Ҡ����K�n-�3�CMKe{>��T�6��IŘ��&�(zI�7z;R;�W1���ΌQո��q�Z�63a�A��‼��e*0��tIn����ֻ��pRcZ�r4����N��J�D
6�jTK��N�
�����^K���0;y�9m9p�LL�e۟
�e*c6�p`]�n1�C��|	e�ݥ@lf�>X�\�=ð���DE���f�Sd�u��d�F\d˙�8p�ڠ>��`U�
�����R�7t�&&�2a�srt`Wgwr�����.R�^�&�H����a�0����]�����b8c��c�8����r9��:0+��%����Nc�	5Zσn	rF�=$���T�l0*�{:0:�unpH�j�@ln��s�n|0;~�T�n�D��(�b!�ܝ���9׾p�V���=@�	H0�
K� � {��o���-�i�����>��T�l0*�丒���߮�̙ͽ�q�e�d8C�[�OjZ��76��q!�D�J&��.5�'/���N��K������GU����k�E�t����Aܝ�����((n�D�Ôq�幊�:0+����J��͆嬡��4����(�����R�N���s��4�L��|pHS����/=��.6ga�W80+����|J�<��� ������d٦�$���  �w��\�2]N)W��UW��rkU�u���yʞ�H]����A����Hy���N��%Kg@q�]M��+����P:�)��ۄ㧕ԏb��]�(W��5���ܗ!Ee�����]86�R۝�l�۬�jW�;Jt���������e�V�\�HI��~}�¢��N��\��p˲Y��\�\�aX�sw��5���+b���k=]΂���}������`Ww)P�ݡʕ
%��.(�
�����S=$꺧�9Ď]ֺ�-�)EI>����J��^C�p`]�����b_C����Ҡ63a�W80�qG�)0=��.f861��E�0*���*��J���-�s�c�D8LG�b�v�����v�޴k`l�g����ȓ��[��+<��Z`W��Gn��Zix��bGr�?��9�h�F@	�G�'Jw��}Ä�WT$�3�G����(��������T��K�p`oq�Tu^�$q��G�Fl0;��ݶ��e*q�T������P��Z���L��*l^C ���ӉR�qA��[�|����s��th������f�ٛ3�-�R�e���0+�����`U�!�w1���8d̾2�;{�%���{��;���.2e���6���W82����we���������H�B!�v 3�{� ��w�9�S� Fp��_� z�D�or3(�Yʀ��9|=	$��"�H1HA���		�ǭ�P�H�x�07N8�F!�,l���	 ��v�1L\h�z�I�%�Á$
$F�X����F@!U���,�F�Oz����끂��k*�(��E� I��$"hE��$=m�q�'B�^��21�BO}�0`H�	� �	���Hz�E�p=�! �9zȑ1� &�h�`v���}����u�"��(r{��T )��?�]" ��@|�}�l����I'�����<��k���Y��v�$��^��|�P���"��1��n��Ƙ]�������\F�7�&{j<�m!÷ �v�p�GG�����Tn����#r�2Ә�m�r���* ��`U��i��[��8�m\�zd�;����o
��J��Ē�/�TC%DL59s@^φe���e* �r��jId��L)��7q�u�9'v�|͓��P�*�"�BBI"����H+$����֨H�"�����ŊF(@ � ���P�	$ �,D�G���y�ٖ��_��n6[s��:I����w\$�^�I� ����X#q �-4��)�K�"s��<�� ��ze��N��17e�df�Ј5@�,
����m0���@xN����3�t��=3� $wl����w�#�� $~�
�!���({Z`V^T�Ǳ��a��ڝD���4����7k�e�hs��8�]�3����I�Ȝ>�w�O6�`�@xx@Do�L@>���R&�T�  �n���*�F��vn��I�&F�i�Ī�6sa��}����vuV�4���vS�eb����)�;Y�GS�D�ݲ7X�s��6:q�tX �=P�۱5�c�m���C������/�Y��&�����U�Zy �7k��x{tI$s��ca'bN���f�
�5z�����m.�7z���hr��� ���\��4��8ѯ,ؠ��.(\�-G�A~�����l̭F�I�jH����v���;��[Z���nq��G�v�m��*y��z.�u��p�dRs,�SͿX;�`��z�~5�5��*��X;��l��/ ��K�����A��lr
�b������N�L �P59n���l�b<϶�����XR��)J��h~G`nȯ��(���n��~����:'Gz�h��H)�{��v��3��[@n���Q.!s�1i��wk��}���P�$A��P�~݃��y��`��K#�p_U�l""[H�QD����n8"�v�r%����\aD'����q�m�"R|/��s3,|��Ն��.�ȹ��`��O7���YW3�T�5��tu��>s�7����'vOP1���߾}<�砹���J �077��;q�Ͼ�~T�f��i9$��}�`�g���Zy����_�&��%�"m3o.v����ݖ��ٸ�̤�u{��B��E����~T�{��X�u�q0�B#���ZynX;�`�lʝf4q��˗`��9�um�A�a�z~^���1�	3xu���;��:���@N�*���_�|�N����	��Y�7n��̭C��1}���١���A)��HN���5�l�{����vEt��Ms�Db��'u��9�ʼy�e��� �F�sE0��`n�n�;r�.]��*}�p��=	n�rF���o�.�%�-�/���xq"�8˰w�O3��;�`�n��"�&3Gش�>�w,�繧�� z����}y�]��Lɶ�Ŵ �>έ�IL)�g
܇l�n���W�"1��KnO1<=(�m���l��53��#b-4���T��=��;�m�N^��܉�<�F�'c-sxr{*�n�ƍ��FÍ�<��W'��1�^�m��T8�B��/H�{C�"�H4f�y�ѮnyΌ��.�"����G�82Φu��2�.��g3�68�U���k�ۺyq\�mנcR8�E�����ܰ����*yޟ��cfڀ�:>۰�`�ʞgٰ���N7�E .�ߕ<�f�߶�>ۧcI��bt}V�w2�߶�3.�n:�a����<�݃�[ ̻2uo��z�w�I4��	�a7$���bzݠ���n���خNz{R���n����o��uw�~rY���[���)IJI�����~~o�����dV��T`$E"
�4AD�<���%���A߿X/��P$����ܖb�x��� ���ܺrQF�*�f��m�~�r���\��sj1�b��s�.���3�O3��>�	: &�V��ݹģ�p���z��N%��q�s�g��3�� .�7�\�sl��wNƒq�PGEŧ��w6�.]��f��P��.]��l���9�s��u1���i�W��]w��34ݩ$�f�<-���P���ޡ`�[$D��R@.]�8�<ϳ`�m�ZsR�ۢKu��@tKݶq�����^%�GFZ�[����
3$踴���;�d<�v�c���NE.]��l��3�O;�~�h�P"�G�vr����hu͚��R����" D�W���y���0@ ����'a)�D1A��ǧ�.A�� �vq�����m�l�m���� <s<��D��z4�	y^�l��P��j �j2�d[�!��`˿�Eŧ�̬�6��6�I�����s����'L_o�X=�QIH&�$c/G>B�O�`�t���*Ae�fN���y�e��k��.�ߕuaq�n(c/���1�h.͘�`���8$�	�Q���� ���A����Q?����"r��?��u�^���<3!��t1��0R,�@��P@��	 �IO$-", �G�
% A H� �2yယ��`�<�5 ���F 6 /G%Sb�$�F"������	  ����!

�(��
� ������b(Qb(� F ����� ���
u \�"d EHE#	2+��:"�Quo��3�X?����� �ȟ@�����<��<A?�Q�~b��V�Ȩ���Q�
7��D���=���x��W�B�5��P��O�?�QW���~vC��`���N�a�����J��
 �^ ��?�_����`����
 �?�Hx� A������?�O�?���?γ������ �~��?�?��������?�"�Q A���?������Ht��*�������#	�K���m?�t�W^s��z�
����O�'T�v������y7�Q�K�
�*$�$��$�²HI""B H	  0��ح�D@Y��@�����	d$@�!	 aI@�dE���I���	�E �EF =�QEUY I$�	!	E$AaAP �Ad@FAU�P$�H@�B0�P!U	 $@FADaT�TD� �XAdHAI@!AA		��DY 		E@Q�DRE	HA�F�(��`(�(�������`�E�T��@ (�P ����� ����"�V(�
,U���� �"�A��D��(����`�`���F�`(�A��Ā�@
�R(�*�D (��"�
� �@(� 
������ 
D �@��AX�,P �D",Q"(0 $X�Fw� �m'_����n��t����~��DP�s0��?g�~�������R��?c���?�_�i����'���_����� �#��P����������7�?�4����{J��?���Q���������2����_��n�$@G�~
(@��'���'�?������ާ��1�ǥ�P
#���D����H���$����O�槇!���_�D@A?u���I*~��N~EDF�!������T	�M��C��p�Ǩ�JG18�!�����#�Α����E��PT��1��?�����ʪ����^�����]���?��O���_���?��aS�?�����A A�� ��?�҈��D?��?{�#����?����/�C�/�����R� d2}�0���6��{��i�?���q���h� ��3����C��������;��ڝ���a�48��s�@���G� �@G���q���޾A�P�w9������p���7�uG��ć�_���B�/��ܑN$3֖�